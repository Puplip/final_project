module gameoverlut (input [23:0] in, input Clk, output out);


always_ff @ (posedge Clk) begin
case (in)

24'h00c01a: out <= 1'b1;
24'h00d01a: out <= 1'b1;
24'h00e01a: out <= 1'b1;
24'h00f01a: out <= 1'b1;
24'h01001a: out <= 1'b1;
24'h01101a: out <= 1'b1;
24'h01201a: out <= 1'b1;
24'h01301a: out <= 1'b1;
24'h01401a: out <= 1'b1;
24'h01501a: out <= 1'b1;
24'h01601a: out <= 1'b1;
24'h01701a: out <= 1'b1;
24'h01801a: out <= 1'b1;
24'h02201a: out <= 1'b1;
24'h02301a: out <= 1'b1;
24'h02401a: out <= 1'b1;
24'h02501a: out <= 1'b1;
24'h02601a: out <= 1'b1;
24'h02701a: out <= 1'b1;
24'h02801a: out <= 1'b1;
24'h02901a: out <= 1'b1;
24'h03201a: out <= 1'b1;
24'h03301a: out <= 1'b1;
24'h03401a: out <= 1'b1;
24'h03501a: out <= 1'b1;
24'h03601a: out <= 1'b1;
24'h03701a: out <= 1'b1;
24'h03f01a: out <= 1'b1;
24'h04001a: out <= 1'b1;
24'h04101a: out <= 1'b1;
24'h04201a: out <= 1'b1;
24'h04301a: out <= 1'b1;
24'h04401a: out <= 1'b1;
24'h04801a: out <= 1'b1;
24'h04901a: out <= 1'b1;
24'h04a01a: out <= 1'b1;
24'h04b01a: out <= 1'b1;
24'h04c01a: out <= 1'b1;
24'h04d01a: out <= 1'b1;
24'h04e01a: out <= 1'b1;
24'h04f01a: out <= 1'b1;
24'h05001a: out <= 1'b1;
24'h05101a: out <= 1'b1;
24'h05201a: out <= 1'b1;
24'h05301a: out <= 1'b1;
24'h05401a: out <= 1'b1;
24'h05501a: out <= 1'b1;
24'h05601a: out <= 1'b1;
24'h05701a: out <= 1'b1;
24'h05801a: out <= 1'b1;
24'h05901a: out <= 1'b1;
24'h05a01a: out <= 1'b1;
24'h00b01b: out <= 1'b1;
24'h00c01b: out <= 1'b1;
24'h00d01b: out <= 1'b1;
24'h00e01b: out <= 1'b1;
24'h00f01b: out <= 1'b1;
24'h01001b: out <= 1'b1;
24'h01101b: out <= 1'b1;
24'h01201b: out <= 1'b1;
24'h01301b: out <= 1'b1;
24'h01401b: out <= 1'b1;
24'h01501b: out <= 1'b1;
24'h01601b: out <= 1'b1;
24'h01701b: out <= 1'b1;
24'h01801b: out <= 1'b1;
24'h01901b: out <= 1'b1;
24'h02101b: out <= 1'b1;
24'h02201b: out <= 1'b1;
24'h02301b: out <= 1'b1;
24'h02401b: out <= 1'b1;
24'h02501b: out <= 1'b1;
24'h02601b: out <= 1'b1;
24'h02701b: out <= 1'b1;
24'h02801b: out <= 1'b1;
24'h02901b: out <= 1'b1;
24'h02a01b: out <= 1'b1;
24'h03201b: out <= 1'b1;
24'h03301b: out <= 1'b1;
24'h03401b: out <= 1'b1;
24'h03501b: out <= 1'b1;
24'h03601b: out <= 1'b1;
24'h03701b: out <= 1'b1;
24'h03801b: out <= 1'b1;
24'h03f01b: out <= 1'b1;
24'h04001b: out <= 1'b1;
24'h04101b: out <= 1'b1;
24'h04201b: out <= 1'b1;
24'h04301b: out <= 1'b1;
24'h04401b: out <= 1'b1;
24'h04501b: out <= 1'b1;
24'h04701b: out <= 1'b1;
24'h04801b: out <= 1'b1;
24'h04901b: out <= 1'b1;
24'h04a01b: out <= 1'b1;
24'h04b01b: out <= 1'b1;
24'h04c01b: out <= 1'b1;
24'h04d01b: out <= 1'b1;
24'h04e01b: out <= 1'b1;
24'h04f01b: out <= 1'b1;
24'h05001b: out <= 1'b1;
24'h05101b: out <= 1'b1;
24'h05201b: out <= 1'b1;
24'h05301b: out <= 1'b1;
24'h05401b: out <= 1'b1;
24'h05501b: out <= 1'b1;
24'h05601b: out <= 1'b1;
24'h05701b: out <= 1'b1;
24'h05801b: out <= 1'b1;
24'h05901b: out <= 1'b1;
24'h05a01b: out <= 1'b1;
24'h05b01b: out <= 1'b1;
24'h00b01c: out <= 1'b1;
24'h00c01c: out <= 1'b1;
24'h00d01c: out <= 1'b1;
24'h00e01c: out <= 1'b1;
24'h00f01c: out <= 1'b1;
24'h01001c: out <= 1'b1;
24'h01101c: out <= 1'b1;
24'h01201c: out <= 1'b1;
24'h01301c: out <= 1'b1;
24'h01401c: out <= 1'b1;
24'h01501c: out <= 1'b1;
24'h01601c: out <= 1'b1;
24'h01701c: out <= 1'b1;
24'h01801c: out <= 1'b1;
24'h01901c: out <= 1'b1;
24'h02101c: out <= 1'b1;
24'h02201c: out <= 1'b1;
24'h02301c: out <= 1'b1;
24'h02401c: out <= 1'b1;
24'h02501c: out <= 1'b1;
24'h02601c: out <= 1'b1;
24'h02701c: out <= 1'b1;
24'h02801c: out <= 1'b1;
24'h02901c: out <= 1'b1;
24'h02a01c: out <= 1'b1;
24'h03201c: out <= 1'b1;
24'h03301c: out <= 1'b1;
24'h03401c: out <= 1'b1;
24'h03501c: out <= 1'b1;
24'h03601c: out <= 1'b1;
24'h03701c: out <= 1'b1;
24'h03801c: out <= 1'b1;
24'h03f01c: out <= 1'b1;
24'h04001c: out <= 1'b1;
24'h04101c: out <= 1'b1;
24'h04201c: out <= 1'b1;
24'h04301c: out <= 1'b1;
24'h04401c: out <= 1'b1;
24'h04501c: out <= 1'b1;
24'h04701c: out <= 1'b1;
24'h04801c: out <= 1'b1;
24'h04901c: out <= 1'b1;
24'h04a01c: out <= 1'b1;
24'h04b01c: out <= 1'b1;
24'h04c01c: out <= 1'b1;
24'h04d01c: out <= 1'b1;
24'h04e01c: out <= 1'b1;
24'h04f01c: out <= 1'b1;
24'h05001c: out <= 1'b1;
24'h05101c: out <= 1'b1;
24'h05201c: out <= 1'b1;
24'h05301c: out <= 1'b1;
24'h05401c: out <= 1'b1;
24'h05501c: out <= 1'b1;
24'h05601c: out <= 1'b1;
24'h05701c: out <= 1'b1;
24'h05801c: out <= 1'b1;
24'h05901c: out <= 1'b1;
24'h05a01c: out <= 1'b1;
24'h05b01c: out <= 1'b1;
24'h00901d: out <= 1'b1;
24'h00a01d: out <= 1'b1;
24'h00b01d: out <= 1'b1;
24'h00c01d: out <= 1'b1;
24'h00d01d: out <= 1'b1;
24'h00e01d: out <= 1'b1;
24'h00f01d: out <= 1'b1;
24'h01001d: out <= 1'b1;
24'h01101d: out <= 1'b1;
24'h01201d: out <= 1'b1;
24'h01301d: out <= 1'b1;
24'h01401d: out <= 1'b1;
24'h01501d: out <= 1'b1;
24'h01601d: out <= 1'b1;
24'h01701d: out <= 1'b1;
24'h01801d: out <= 1'b1;
24'h01901d: out <= 1'b1;
24'h01f01d: out <= 1'b1;
24'h02001d: out <= 1'b1;
24'h02101d: out <= 1'b1;
24'h02201d: out <= 1'b1;
24'h02301d: out <= 1'b1;
24'h02401d: out <= 1'b1;
24'h02501d: out <= 1'b1;
24'h02601d: out <= 1'b1;
24'h02701d: out <= 1'b1;
24'h02801d: out <= 1'b1;
24'h02901d: out <= 1'b1;
24'h02a01d: out <= 1'b1;
24'h02b01d: out <= 1'b1;
24'h02c01d: out <= 1'b1;
24'h03201d: out <= 1'b1;
24'h03301d: out <= 1'b1;
24'h03401d: out <= 1'b1;
24'h03501d: out <= 1'b1;
24'h03601d: out <= 1'b1;
24'h03701d: out <= 1'b1;
24'h03801d: out <= 1'b1;
24'h03901d: out <= 1'b1;
24'h03a01d: out <= 1'b1;
24'h03c01d: out <= 1'b1;
24'h03d01d: out <= 1'b1;
24'h03e01d: out <= 1'b1;
24'h03f01d: out <= 1'b1;
24'h04001d: out <= 1'b1;
24'h04101d: out <= 1'b1;
24'h04201d: out <= 1'b1;
24'h04301d: out <= 1'b1;
24'h04401d: out <= 1'b1;
24'h04501d: out <= 1'b1;
24'h04701d: out <= 1'b1;
24'h04801d: out <= 1'b1;
24'h04901d: out <= 1'b1;
24'h04a01d: out <= 1'b1;
24'h04b01d: out <= 1'b1;
24'h04c01d: out <= 1'b1;
24'h04d01d: out <= 1'b1;
24'h04e01d: out <= 1'b1;
24'h04f01d: out <= 1'b1;
24'h05001d: out <= 1'b1;
24'h05101d: out <= 1'b1;
24'h05201d: out <= 1'b1;
24'h05301d: out <= 1'b1;
24'h05401d: out <= 1'b1;
24'h05501d: out <= 1'b1;
24'h05601d: out <= 1'b1;
24'h05701d: out <= 1'b1;
24'h05801d: out <= 1'b1;
24'h05901d: out <= 1'b1;
24'h05a01d: out <= 1'b1;
24'h05b01d: out <= 1'b1;
24'h00801e: out <= 1'b1;
24'h00901e: out <= 1'b1;
24'h00a01e: out <= 1'b1;
24'h00b01e: out <= 1'b1;
24'h00c01e: out <= 1'b1;
24'h00d01e: out <= 1'b1;
24'h00e01e: out <= 1'b1;
24'h00f01e: out <= 1'b1;
24'h01001e: out <= 1'b1;
24'h01101e: out <= 1'b1;
24'h01201e: out <= 1'b1;
24'h01301e: out <= 1'b1;
24'h01401e: out <= 1'b1;
24'h01501e: out <= 1'b1;
24'h01601e: out <= 1'b1;
24'h01701e: out <= 1'b1;
24'h01801e: out <= 1'b1;
24'h01901e: out <= 1'b1;
24'h01e01e: out <= 1'b1;
24'h01f01e: out <= 1'b1;
24'h02001e: out <= 1'b1;
24'h02101e: out <= 1'b1;
24'h02201e: out <= 1'b1;
24'h02301e: out <= 1'b1;
24'h02401e: out <= 1'b1;
24'h02501e: out <= 1'b1;
24'h02601e: out <= 1'b1;
24'h02701e: out <= 1'b1;
24'h02801e: out <= 1'b1;
24'h02901e: out <= 1'b1;
24'h02a01e: out <= 1'b1;
24'h02b01e: out <= 1'b1;
24'h02c01e: out <= 1'b1;
24'h03201e: out <= 1'b1;
24'h03301e: out <= 1'b1;
24'h03401e: out <= 1'b1;
24'h03501e: out <= 1'b1;
24'h03601e: out <= 1'b1;
24'h03701e: out <= 1'b1;
24'h03801e: out <= 1'b1;
24'h03901e: out <= 1'b1;
24'h03a01e: out <= 1'b1;
24'h03c01e: out <= 1'b1;
24'h03d01e: out <= 1'b1;
24'h03e01e: out <= 1'b1;
24'h03f01e: out <= 1'b1;
24'h04001e: out <= 1'b1;
24'h04101e: out <= 1'b1;
24'h04201e: out <= 1'b1;
24'h04301e: out <= 1'b1;
24'h04401e: out <= 1'b1;
24'h04501e: out <= 1'b1;
24'h04701e: out <= 1'b1;
24'h04801e: out <= 1'b1;
24'h04901e: out <= 1'b1;
24'h04a01e: out <= 1'b1;
24'h04b01e: out <= 1'b1;
24'h04c01e: out <= 1'b1;
24'h04d01e: out <= 1'b1;
24'h04e01e: out <= 1'b1;
24'h04f01e: out <= 1'b1;
24'h05001e: out <= 1'b1;
24'h05101e: out <= 1'b1;
24'h05201e: out <= 1'b1;
24'h05301e: out <= 1'b1;
24'h05401e: out <= 1'b1;
24'h05501e: out <= 1'b1;
24'h05601e: out <= 1'b1;
24'h05701e: out <= 1'b1;
24'h05801e: out <= 1'b1;
24'h05901e: out <= 1'b1;
24'h05a01e: out <= 1'b1;
24'h00801f: out <= 1'b1;
24'h00901f: out <= 1'b1;
24'h00a01f: out <= 1'b1;
24'h00b01f: out <= 1'b1;
24'h00c01f: out <= 1'b1;
24'h00d01f: out <= 1'b1;
24'h00e01f: out <= 1'b1;
24'h00f01f: out <= 1'b1;
24'h01e01f: out <= 1'b1;
24'h01f01f: out <= 1'b1;
24'h02001f: out <= 1'b1;
24'h02101f: out <= 1'b1;
24'h02201f: out <= 1'b1;
24'h02301f: out <= 1'b1;
24'h02401f: out <= 1'b1;
24'h02601f: out <= 1'b1;
24'h02701f: out <= 1'b1;
24'h02801f: out <= 1'b1;
24'h02901f: out <= 1'b1;
24'h02a01f: out <= 1'b1;
24'h02b01f: out <= 1'b1;
24'h02c01f: out <= 1'b1;
24'h03201f: out <= 1'b1;
24'h03301f: out <= 1'b1;
24'h03401f: out <= 1'b1;
24'h03501f: out <= 1'b1;
24'h03601f: out <= 1'b1;
24'h03701f: out <= 1'b1;
24'h03801f: out <= 1'b1;
24'h03901f: out <= 1'b1;
24'h03a01f: out <= 1'b1;
24'h03c01f: out <= 1'b1;
24'h03d01f: out <= 1'b1;
24'h03e01f: out <= 1'b1;
24'h03f01f: out <= 1'b1;
24'h04001f: out <= 1'b1;
24'h04101f: out <= 1'b1;
24'h04201f: out <= 1'b1;
24'h04301f: out <= 1'b1;
24'h04401f: out <= 1'b1;
24'h04501f: out <= 1'b1;
24'h04701f: out <= 1'b1;
24'h04801f: out <= 1'b1;
24'h04901f: out <= 1'b1;
24'h04a01f: out <= 1'b1;
24'h04b01f: out <= 1'b1;
24'h04c01f: out <= 1'b1;
24'h04d01f: out <= 1'b1;
24'h04e01f: out <= 1'b1;
24'h006020: out <= 1'b1;
24'h007020: out <= 1'b1;
24'h008020: out <= 1'b1;
24'h009020: out <= 1'b1;
24'h00a020: out <= 1'b1;
24'h00b020: out <= 1'b1;
24'h00c020: out <= 1'b1;
24'h00d020: out <= 1'b1;
24'h00e020: out <= 1'b1;
24'h01c020: out <= 1'b1;
24'h01d020: out <= 1'b1;
24'h01e020: out <= 1'b1;
24'h01f020: out <= 1'b1;
24'h020020: out <= 1'b1;
24'h021020: out <= 1'b1;
24'h022020: out <= 1'b1;
24'h023020: out <= 1'b1;
24'h024020: out <= 1'b1;
24'h026020: out <= 1'b1;
24'h027020: out <= 1'b1;
24'h028020: out <= 1'b1;
24'h029020: out <= 1'b1;
24'h02a020: out <= 1'b1;
24'h02b020: out <= 1'b1;
24'h02c020: out <= 1'b1;
24'h02d020: out <= 1'b1;
24'h02e020: out <= 1'b1;
24'h02f020: out <= 1'b1;
24'h032020: out <= 1'b1;
24'h033020: out <= 1'b1;
24'h034020: out <= 1'b1;
24'h035020: out <= 1'b1;
24'h036020: out <= 1'b1;
24'h037020: out <= 1'b1;
24'h038020: out <= 1'b1;
24'h039020: out <= 1'b1;
24'h03a020: out <= 1'b1;
24'h03b020: out <= 1'b1;
24'h03c020: out <= 1'b1;
24'h03d020: out <= 1'b1;
24'h03e020: out <= 1'b1;
24'h03f020: out <= 1'b1;
24'h040020: out <= 1'b1;
24'h041020: out <= 1'b1;
24'h042020: out <= 1'b1;
24'h043020: out <= 1'b1;
24'h044020: out <= 1'b1;
24'h045020: out <= 1'b1;
24'h047020: out <= 1'b1;
24'h048020: out <= 1'b1;
24'h049020: out <= 1'b1;
24'h04a020: out <= 1'b1;
24'h04b020: out <= 1'b1;
24'h04c020: out <= 1'b1;
24'h04d020: out <= 1'b1;
24'h04e020: out <= 1'b1;
24'h006021: out <= 1'b1;
24'h007021: out <= 1'b1;
24'h008021: out <= 1'b1;
24'h009021: out <= 1'b1;
24'h00a021: out <= 1'b1;
24'h00b021: out <= 1'b1;
24'h00c021: out <= 1'b1;
24'h01c021: out <= 1'b1;
24'h01d021: out <= 1'b1;
24'h01e021: out <= 1'b1;
24'h01f021: out <= 1'b1;
24'h020021: out <= 1'b1;
24'h021021: out <= 1'b1;
24'h022021: out <= 1'b1;
24'h029021: out <= 1'b1;
24'h02a021: out <= 1'b1;
24'h02b021: out <= 1'b1;
24'h02c021: out <= 1'b1;
24'h02d021: out <= 1'b1;
24'h02e021: out <= 1'b1;
24'h02f021: out <= 1'b1;
24'h032021: out <= 1'b1;
24'h033021: out <= 1'b1;
24'h034021: out <= 1'b1;
24'h035021: out <= 1'b1;
24'h036021: out <= 1'b1;
24'h037021: out <= 1'b1;
24'h038021: out <= 1'b1;
24'h039021: out <= 1'b1;
24'h03a021: out <= 1'b1;
24'h03b021: out <= 1'b1;
24'h03c021: out <= 1'b1;
24'h03d021: out <= 1'b1;
24'h03e021: out <= 1'b1;
24'h03f021: out <= 1'b1;
24'h040021: out <= 1'b1;
24'h041021: out <= 1'b1;
24'h042021: out <= 1'b1;
24'h043021: out <= 1'b1;
24'h044021: out <= 1'b1;
24'h045021: out <= 1'b1;
24'h047021: out <= 1'b1;
24'h048021: out <= 1'b1;
24'h049021: out <= 1'b1;
24'h04a021: out <= 1'b1;
24'h04b021: out <= 1'b1;
24'h04c021: out <= 1'b1;
24'h04d021: out <= 1'b1;
24'h04e021: out <= 1'b1;
24'h006022: out <= 1'b1;
24'h007022: out <= 1'b1;
24'h008022: out <= 1'b1;
24'h009022: out <= 1'b1;
24'h00a022: out <= 1'b1;
24'h00b022: out <= 1'b1;
24'h00c022: out <= 1'b1;
24'h011022: out <= 1'b1;
24'h012022: out <= 1'b1;
24'h013022: out <= 1'b1;
24'h014022: out <= 1'b1;
24'h015022: out <= 1'b1;
24'h016022: out <= 1'b1;
24'h017022: out <= 1'b1;
24'h018022: out <= 1'b1;
24'h019022: out <= 1'b1;
24'h01c022: out <= 1'b1;
24'h01d022: out <= 1'b1;
24'h01e022: out <= 1'b1;
24'h01f022: out <= 1'b1;
24'h020022: out <= 1'b1;
24'h021022: out <= 1'b1;
24'h022022: out <= 1'b1;
24'h029022: out <= 1'b1;
24'h02a022: out <= 1'b1;
24'h02b022: out <= 1'b1;
24'h02c022: out <= 1'b1;
24'h02d022: out <= 1'b1;
24'h02e022: out <= 1'b1;
24'h02f022: out <= 1'b1;
24'h032022: out <= 1'b1;
24'h033022: out <= 1'b1;
24'h034022: out <= 1'b1;
24'h035022: out <= 1'b1;
24'h036022: out <= 1'b1;
24'h037022: out <= 1'b1;
24'h038022: out <= 1'b1;
24'h039022: out <= 1'b1;
24'h03a022: out <= 1'b1;
24'h03b022: out <= 1'b1;
24'h03c022: out <= 1'b1;
24'h03d022: out <= 1'b1;
24'h03e022: out <= 1'b1;
24'h03f022: out <= 1'b1;
24'h040022: out <= 1'b1;
24'h041022: out <= 1'b1;
24'h042022: out <= 1'b1;
24'h043022: out <= 1'b1;
24'h044022: out <= 1'b1;
24'h045022: out <= 1'b1;
24'h047022: out <= 1'b1;
24'h048022: out <= 1'b1;
24'h049022: out <= 1'b1;
24'h04a022: out <= 1'b1;
24'h04b022: out <= 1'b1;
24'h04c022: out <= 1'b1;
24'h04d022: out <= 1'b1;
24'h04e022: out <= 1'b1;
24'h04f022: out <= 1'b1;
24'h050022: out <= 1'b1;
24'h051022: out <= 1'b1;
24'h052022: out <= 1'b1;
24'h053022: out <= 1'b1;
24'h054022: out <= 1'b1;
24'h055022: out <= 1'b1;
24'h056022: out <= 1'b1;
24'h057022: out <= 1'b1;
24'h058022: out <= 1'b1;
24'h006023: out <= 1'b1;
24'h007023: out <= 1'b1;
24'h008023: out <= 1'b1;
24'h009023: out <= 1'b1;
24'h00a023: out <= 1'b1;
24'h00b023: out <= 1'b1;
24'h00c023: out <= 1'b1;
24'h010023: out <= 1'b1;
24'h011023: out <= 1'b1;
24'h012023: out <= 1'b1;
24'h013023: out <= 1'b1;
24'h014023: out <= 1'b1;
24'h015023: out <= 1'b1;
24'h016023: out <= 1'b1;
24'h017023: out <= 1'b1;
24'h018023: out <= 1'b1;
24'h019023: out <= 1'b1;
24'h01c023: out <= 1'b1;
24'h01d023: out <= 1'b1;
24'h01e023: out <= 1'b1;
24'h01f023: out <= 1'b1;
24'h020023: out <= 1'b1;
24'h021023: out <= 1'b1;
24'h022023: out <= 1'b1;
24'h029023: out <= 1'b1;
24'h02a023: out <= 1'b1;
24'h02b023: out <= 1'b1;
24'h02c023: out <= 1'b1;
24'h02d023: out <= 1'b1;
24'h02e023: out <= 1'b1;
24'h02f023: out <= 1'b1;
24'h032023: out <= 1'b1;
24'h033023: out <= 1'b1;
24'h034023: out <= 1'b1;
24'h035023: out <= 1'b1;
24'h036023: out <= 1'b1;
24'h037023: out <= 1'b1;
24'h038023: out <= 1'b1;
24'h039023: out <= 1'b1;
24'h03a023: out <= 1'b1;
24'h03b023: out <= 1'b1;
24'h03c023: out <= 1'b1;
24'h03d023: out <= 1'b1;
24'h03e023: out <= 1'b1;
24'h03f023: out <= 1'b1;
24'h040023: out <= 1'b1;
24'h041023: out <= 1'b1;
24'h042023: out <= 1'b1;
24'h043023: out <= 1'b1;
24'h044023: out <= 1'b1;
24'h045023: out <= 1'b1;
24'h047023: out <= 1'b1;
24'h048023: out <= 1'b1;
24'h049023: out <= 1'b1;
24'h04a023: out <= 1'b1;
24'h04b023: out <= 1'b1;
24'h04c023: out <= 1'b1;
24'h04d023: out <= 1'b1;
24'h04e023: out <= 1'b1;
24'h04f023: out <= 1'b1;
24'h050023: out <= 1'b1;
24'h051023: out <= 1'b1;
24'h052023: out <= 1'b1;
24'h053023: out <= 1'b1;
24'h054023: out <= 1'b1;
24'h055023: out <= 1'b1;
24'h056023: out <= 1'b1;
24'h057023: out <= 1'b1;
24'h058023: out <= 1'b1;
24'h006024: out <= 1'b1;
24'h007024: out <= 1'b1;
24'h008024: out <= 1'b1;
24'h009024: out <= 1'b1;
24'h00a024: out <= 1'b1;
24'h00b024: out <= 1'b1;
24'h00c024: out <= 1'b1;
24'h010024: out <= 1'b1;
24'h011024: out <= 1'b1;
24'h012024: out <= 1'b1;
24'h013024: out <= 1'b1;
24'h014024: out <= 1'b1;
24'h015024: out <= 1'b1;
24'h016024: out <= 1'b1;
24'h017024: out <= 1'b1;
24'h018024: out <= 1'b1;
24'h019024: out <= 1'b1;
24'h01c024: out <= 1'b1;
24'h01d024: out <= 1'b1;
24'h01e024: out <= 1'b1;
24'h01f024: out <= 1'b1;
24'h020024: out <= 1'b1;
24'h021024: out <= 1'b1;
24'h022024: out <= 1'b1;
24'h029024: out <= 1'b1;
24'h02a024: out <= 1'b1;
24'h02b024: out <= 1'b1;
24'h02c024: out <= 1'b1;
24'h02d024: out <= 1'b1;
24'h02e024: out <= 1'b1;
24'h02f024: out <= 1'b1;
24'h032024: out <= 1'b1;
24'h033024: out <= 1'b1;
24'h034024: out <= 1'b1;
24'h035024: out <= 1'b1;
24'h036024: out <= 1'b1;
24'h037024: out <= 1'b1;
24'h038024: out <= 1'b1;
24'h039024: out <= 1'b1;
24'h03a024: out <= 1'b1;
24'h03b024: out <= 1'b1;
24'h03c024: out <= 1'b1;
24'h03d024: out <= 1'b1;
24'h03e024: out <= 1'b1;
24'h03f024: out <= 1'b1;
24'h040024: out <= 1'b1;
24'h041024: out <= 1'b1;
24'h042024: out <= 1'b1;
24'h043024: out <= 1'b1;
24'h044024: out <= 1'b1;
24'h045024: out <= 1'b1;
24'h047024: out <= 1'b1;
24'h048024: out <= 1'b1;
24'h049024: out <= 1'b1;
24'h04a024: out <= 1'b1;
24'h04b024: out <= 1'b1;
24'h04c024: out <= 1'b1;
24'h04d024: out <= 1'b1;
24'h04e024: out <= 1'b1;
24'h04f024: out <= 1'b1;
24'h050024: out <= 1'b1;
24'h051024: out <= 1'b1;
24'h052024: out <= 1'b1;
24'h053024: out <= 1'b1;
24'h054024: out <= 1'b1;
24'h055024: out <= 1'b1;
24'h056024: out <= 1'b1;
24'h057024: out <= 1'b1;
24'h058024: out <= 1'b1;
24'h006025: out <= 1'b1;
24'h007025: out <= 1'b1;
24'h008025: out <= 1'b1;
24'h009025: out <= 1'b1;
24'h00a025: out <= 1'b1;
24'h00b025: out <= 1'b1;
24'h00c025: out <= 1'b1;
24'h010025: out <= 1'b1;
24'h011025: out <= 1'b1;
24'h012025: out <= 1'b1;
24'h013025: out <= 1'b1;
24'h014025: out <= 1'b1;
24'h015025: out <= 1'b1;
24'h016025: out <= 1'b1;
24'h017025: out <= 1'b1;
24'h018025: out <= 1'b1;
24'h019025: out <= 1'b1;
24'h01c025: out <= 1'b1;
24'h01d025: out <= 1'b1;
24'h01e025: out <= 1'b1;
24'h01f025: out <= 1'b1;
24'h020025: out <= 1'b1;
24'h021025: out <= 1'b1;
24'h022025: out <= 1'b1;
24'h023025: out <= 1'b1;
24'h024025: out <= 1'b1;
24'h025025: out <= 1'b1;
24'h026025: out <= 1'b1;
24'h027025: out <= 1'b1;
24'h028025: out <= 1'b1;
24'h029025: out <= 1'b1;
24'h02a025: out <= 1'b1;
24'h02b025: out <= 1'b1;
24'h02c025: out <= 1'b1;
24'h02d025: out <= 1'b1;
24'h02e025: out <= 1'b1;
24'h02f025: out <= 1'b1;
24'h032025: out <= 1'b1;
24'h033025: out <= 1'b1;
24'h034025: out <= 1'b1;
24'h035025: out <= 1'b1;
24'h036025: out <= 1'b1;
24'h037025: out <= 1'b1;
24'h038025: out <= 1'b1;
24'h039025: out <= 1'b1;
24'h03a025: out <= 1'b1;
24'h03b025: out <= 1'b1;
24'h03c025: out <= 1'b1;
24'h03d025: out <= 1'b1;
24'h03e025: out <= 1'b1;
24'h03f025: out <= 1'b1;
24'h040025: out <= 1'b1;
24'h041025: out <= 1'b1;
24'h042025: out <= 1'b1;
24'h043025: out <= 1'b1;
24'h044025: out <= 1'b1;
24'h045025: out <= 1'b1;
24'h047025: out <= 1'b1;
24'h048025: out <= 1'b1;
24'h049025: out <= 1'b1;
24'h04a025: out <= 1'b1;
24'h04b025: out <= 1'b1;
24'h04c025: out <= 1'b1;
24'h04d025: out <= 1'b1;
24'h04e025: out <= 1'b1;
24'h04f025: out <= 1'b1;
24'h050025: out <= 1'b1;
24'h051025: out <= 1'b1;
24'h052025: out <= 1'b1;
24'h053025: out <= 1'b1;
24'h054025: out <= 1'b1;
24'h055025: out <= 1'b1;
24'h056025: out <= 1'b1;
24'h057025: out <= 1'b1;
24'h058025: out <= 1'b1;
24'h006026: out <= 1'b1;
24'h007026: out <= 1'b1;
24'h008026: out <= 1'b1;
24'h009026: out <= 1'b1;
24'h00a026: out <= 1'b1;
24'h00b026: out <= 1'b1;
24'h00c026: out <= 1'b1;
24'h011026: out <= 1'b1;
24'h012026: out <= 1'b1;
24'h013026: out <= 1'b1;
24'h014026: out <= 1'b1;
24'h015026: out <= 1'b1;
24'h016026: out <= 1'b1;
24'h017026: out <= 1'b1;
24'h018026: out <= 1'b1;
24'h019026: out <= 1'b1;
24'h01c026: out <= 1'b1;
24'h01d026: out <= 1'b1;
24'h01e026: out <= 1'b1;
24'h01f026: out <= 1'b1;
24'h020026: out <= 1'b1;
24'h021026: out <= 1'b1;
24'h022026: out <= 1'b1;
24'h023026: out <= 1'b1;
24'h024026: out <= 1'b1;
24'h025026: out <= 1'b1;
24'h026026: out <= 1'b1;
24'h027026: out <= 1'b1;
24'h028026: out <= 1'b1;
24'h029026: out <= 1'b1;
24'h02a026: out <= 1'b1;
24'h02b026: out <= 1'b1;
24'h02c026: out <= 1'b1;
24'h02d026: out <= 1'b1;
24'h02e026: out <= 1'b1;
24'h02f026: out <= 1'b1;
24'h032026: out <= 1'b1;
24'h033026: out <= 1'b1;
24'h034026: out <= 1'b1;
24'h035026: out <= 1'b1;
24'h036026: out <= 1'b1;
24'h037026: out <= 1'b1;
24'h038026: out <= 1'b1;
24'h039026: out <= 1'b1;
24'h03a026: out <= 1'b1;
24'h03b026: out <= 1'b1;
24'h03c026: out <= 1'b1;
24'h03d026: out <= 1'b1;
24'h03e026: out <= 1'b1;
24'h03f026: out <= 1'b1;
24'h040026: out <= 1'b1;
24'h041026: out <= 1'b1;
24'h042026: out <= 1'b1;
24'h043026: out <= 1'b1;
24'h044026: out <= 1'b1;
24'h045026: out <= 1'b1;
24'h047026: out <= 1'b1;
24'h048026: out <= 1'b1;
24'h049026: out <= 1'b1;
24'h04a026: out <= 1'b1;
24'h04b026: out <= 1'b1;
24'h04c026: out <= 1'b1;
24'h04d026: out <= 1'b1;
24'h04e026: out <= 1'b1;
24'h04f026: out <= 1'b1;
24'h050026: out <= 1'b1;
24'h051026: out <= 1'b1;
24'h052026: out <= 1'b1;
24'h053026: out <= 1'b1;
24'h054026: out <= 1'b1;
24'h055026: out <= 1'b1;
24'h056026: out <= 1'b1;
24'h057026: out <= 1'b1;
24'h058026: out <= 1'b1;
24'h006027: out <= 1'b1;
24'h007027: out <= 1'b1;
24'h008027: out <= 1'b1;
24'h009027: out <= 1'b1;
24'h00a027: out <= 1'b1;
24'h00b027: out <= 1'b1;
24'h00c027: out <= 1'b1;
24'h013027: out <= 1'b1;
24'h014027: out <= 1'b1;
24'h015027: out <= 1'b1;
24'h016027: out <= 1'b1;
24'h017027: out <= 1'b1;
24'h018027: out <= 1'b1;
24'h019027: out <= 1'b1;
24'h01c027: out <= 1'b1;
24'h01d027: out <= 1'b1;
24'h01e027: out <= 1'b1;
24'h01f027: out <= 1'b1;
24'h020027: out <= 1'b1;
24'h021027: out <= 1'b1;
24'h022027: out <= 1'b1;
24'h023027: out <= 1'b1;
24'h024027: out <= 1'b1;
24'h025027: out <= 1'b1;
24'h026027: out <= 1'b1;
24'h027027: out <= 1'b1;
24'h028027: out <= 1'b1;
24'h029027: out <= 1'b1;
24'h02a027: out <= 1'b1;
24'h02b027: out <= 1'b1;
24'h02c027: out <= 1'b1;
24'h02d027: out <= 1'b1;
24'h02e027: out <= 1'b1;
24'h02f027: out <= 1'b1;
24'h032027: out <= 1'b1;
24'h033027: out <= 1'b1;
24'h034027: out <= 1'b1;
24'h035027: out <= 1'b1;
24'h036027: out <= 1'b1;
24'h037027: out <= 1'b1;
24'h038027: out <= 1'b1;
24'h03a027: out <= 1'b1;
24'h03b027: out <= 1'b1;
24'h03c027: out <= 1'b1;
24'h03d027: out <= 1'b1;
24'h03f027: out <= 1'b1;
24'h040027: out <= 1'b1;
24'h041027: out <= 1'b1;
24'h042027: out <= 1'b1;
24'h043027: out <= 1'b1;
24'h044027: out <= 1'b1;
24'h045027: out <= 1'b1;
24'h047027: out <= 1'b1;
24'h048027: out <= 1'b1;
24'h049027: out <= 1'b1;
24'h04a027: out <= 1'b1;
24'h04b027: out <= 1'b1;
24'h04c027: out <= 1'b1;
24'h04d027: out <= 1'b1;
24'h04e027: out <= 1'b1;
24'h006028: out <= 1'b1;
24'h007028: out <= 1'b1;
24'h008028: out <= 1'b1;
24'h009028: out <= 1'b1;
24'h00a028: out <= 1'b1;
24'h00b028: out <= 1'b1;
24'h00c028: out <= 1'b1;
24'h00d028: out <= 1'b1;
24'h00e028: out <= 1'b1;
24'h013028: out <= 1'b1;
24'h014028: out <= 1'b1;
24'h015028: out <= 1'b1;
24'h016028: out <= 1'b1;
24'h017028: out <= 1'b1;
24'h018028: out <= 1'b1;
24'h019028: out <= 1'b1;
24'h01c028: out <= 1'b1;
24'h01d028: out <= 1'b1;
24'h01e028: out <= 1'b1;
24'h01f028: out <= 1'b1;
24'h020028: out <= 1'b1;
24'h021028: out <= 1'b1;
24'h022028: out <= 1'b1;
24'h023028: out <= 1'b1;
24'h024028: out <= 1'b1;
24'h025028: out <= 1'b1;
24'h026028: out <= 1'b1;
24'h027028: out <= 1'b1;
24'h028028: out <= 1'b1;
24'h029028: out <= 1'b1;
24'h02a028: out <= 1'b1;
24'h02b028: out <= 1'b1;
24'h02c028: out <= 1'b1;
24'h02d028: out <= 1'b1;
24'h02e028: out <= 1'b1;
24'h02f028: out <= 1'b1;
24'h032028: out <= 1'b1;
24'h033028: out <= 1'b1;
24'h034028: out <= 1'b1;
24'h035028: out <= 1'b1;
24'h036028: out <= 1'b1;
24'h037028: out <= 1'b1;
24'h038028: out <= 1'b1;
24'h03a028: out <= 1'b1;
24'h03b028: out <= 1'b1;
24'h03c028: out <= 1'b1;
24'h03d028: out <= 1'b1;
24'h03f028: out <= 1'b1;
24'h040028: out <= 1'b1;
24'h041028: out <= 1'b1;
24'h042028: out <= 1'b1;
24'h043028: out <= 1'b1;
24'h044028: out <= 1'b1;
24'h045028: out <= 1'b1;
24'h047028: out <= 1'b1;
24'h048028: out <= 1'b1;
24'h049028: out <= 1'b1;
24'h04a028: out <= 1'b1;
24'h04b028: out <= 1'b1;
24'h04c028: out <= 1'b1;
24'h04d028: out <= 1'b1;
24'h04e028: out <= 1'b1;
24'h008029: out <= 1'b1;
24'h009029: out <= 1'b1;
24'h00a029: out <= 1'b1;
24'h00b029: out <= 1'b1;
24'h00c029: out <= 1'b1;
24'h00d029: out <= 1'b1;
24'h00e029: out <= 1'b1;
24'h00f029: out <= 1'b1;
24'h013029: out <= 1'b1;
24'h014029: out <= 1'b1;
24'h015029: out <= 1'b1;
24'h016029: out <= 1'b1;
24'h017029: out <= 1'b1;
24'h018029: out <= 1'b1;
24'h019029: out <= 1'b1;
24'h01c029: out <= 1'b1;
24'h01d029: out <= 1'b1;
24'h01e029: out <= 1'b1;
24'h01f029: out <= 1'b1;
24'h020029: out <= 1'b1;
24'h021029: out <= 1'b1;
24'h022029: out <= 1'b1;
24'h029029: out <= 1'b1;
24'h02a029: out <= 1'b1;
24'h02b029: out <= 1'b1;
24'h02c029: out <= 1'b1;
24'h02d029: out <= 1'b1;
24'h02e029: out <= 1'b1;
24'h02f029: out <= 1'b1;
24'h032029: out <= 1'b1;
24'h033029: out <= 1'b1;
24'h034029: out <= 1'b1;
24'h035029: out <= 1'b1;
24'h036029: out <= 1'b1;
24'h037029: out <= 1'b1;
24'h038029: out <= 1'b1;
24'h03f029: out <= 1'b1;
24'h040029: out <= 1'b1;
24'h041029: out <= 1'b1;
24'h042029: out <= 1'b1;
24'h043029: out <= 1'b1;
24'h044029: out <= 1'b1;
24'h045029: out <= 1'b1;
24'h047029: out <= 1'b1;
24'h048029: out <= 1'b1;
24'h049029: out <= 1'b1;
24'h04a029: out <= 1'b1;
24'h04b029: out <= 1'b1;
24'h04c029: out <= 1'b1;
24'h04d029: out <= 1'b1;
24'h04e029: out <= 1'b1;
24'h00802a: out <= 1'b1;
24'h00902a: out <= 1'b1;
24'h00a02a: out <= 1'b1;
24'h00b02a: out <= 1'b1;
24'h00c02a: out <= 1'b1;
24'h00d02a: out <= 1'b1;
24'h00e02a: out <= 1'b1;
24'h00f02a: out <= 1'b1;
24'h01002a: out <= 1'b1;
24'h01102a: out <= 1'b1;
24'h01202a: out <= 1'b1;
24'h01302a: out <= 1'b1;
24'h01402a: out <= 1'b1;
24'h01502a: out <= 1'b1;
24'h01602a: out <= 1'b1;
24'h01702a: out <= 1'b1;
24'h01802a: out <= 1'b1;
24'h01902a: out <= 1'b1;
24'h01c02a: out <= 1'b1;
24'h01d02a: out <= 1'b1;
24'h01e02a: out <= 1'b1;
24'h01f02a: out <= 1'b1;
24'h02002a: out <= 1'b1;
24'h02102a: out <= 1'b1;
24'h02202a: out <= 1'b1;
24'h02902a: out <= 1'b1;
24'h02a02a: out <= 1'b1;
24'h02b02a: out <= 1'b1;
24'h02c02a: out <= 1'b1;
24'h02d02a: out <= 1'b1;
24'h02e02a: out <= 1'b1;
24'h02f02a: out <= 1'b1;
24'h03202a: out <= 1'b1;
24'h03302a: out <= 1'b1;
24'h03402a: out <= 1'b1;
24'h03502a: out <= 1'b1;
24'h03602a: out <= 1'b1;
24'h03702a: out <= 1'b1;
24'h03802a: out <= 1'b1;
24'h03f02a: out <= 1'b1;
24'h04002a: out <= 1'b1;
24'h04102a: out <= 1'b1;
24'h04202a: out <= 1'b1;
24'h04302a: out <= 1'b1;
24'h04402a: out <= 1'b1;
24'h04502a: out <= 1'b1;
24'h04702a: out <= 1'b1;
24'h04802a: out <= 1'b1;
24'h04902a: out <= 1'b1;
24'h04a02a: out <= 1'b1;
24'h04b02a: out <= 1'b1;
24'h04c02a: out <= 1'b1;
24'h04d02a: out <= 1'b1;
24'h04e02a: out <= 1'b1;
24'h04f02a: out <= 1'b1;
24'h05002a: out <= 1'b1;
24'h05102a: out <= 1'b1;
24'h05202a: out <= 1'b1;
24'h05302a: out <= 1'b1;
24'h05402a: out <= 1'b1;
24'h05502a: out <= 1'b1;
24'h05602a: out <= 1'b1;
24'h05702a: out <= 1'b1;
24'h05802a: out <= 1'b1;
24'h05902a: out <= 1'b1;
24'h05a02a: out <= 1'b1;
24'h00902b: out <= 1'b1;
24'h00a02b: out <= 1'b1;
24'h00b02b: out <= 1'b1;
24'h00c02b: out <= 1'b1;
24'h00d02b: out <= 1'b1;
24'h00e02b: out <= 1'b1;
24'h00f02b: out <= 1'b1;
24'h01002b: out <= 1'b1;
24'h01102b: out <= 1'b1;
24'h01202b: out <= 1'b1;
24'h01302b: out <= 1'b1;
24'h01402b: out <= 1'b1;
24'h01502b: out <= 1'b1;
24'h01602b: out <= 1'b1;
24'h01702b: out <= 1'b1;
24'h01802b: out <= 1'b1;
24'h01902b: out <= 1'b1;
24'h01c02b: out <= 1'b1;
24'h01d02b: out <= 1'b1;
24'h01e02b: out <= 1'b1;
24'h01f02b: out <= 1'b1;
24'h02002b: out <= 1'b1;
24'h02102b: out <= 1'b1;
24'h02202b: out <= 1'b1;
24'h02902b: out <= 1'b1;
24'h02a02b: out <= 1'b1;
24'h02b02b: out <= 1'b1;
24'h02c02b: out <= 1'b1;
24'h02d02b: out <= 1'b1;
24'h02e02b: out <= 1'b1;
24'h02f02b: out <= 1'b1;
24'h03202b: out <= 1'b1;
24'h03302b: out <= 1'b1;
24'h03402b: out <= 1'b1;
24'h03502b: out <= 1'b1;
24'h03602b: out <= 1'b1;
24'h03702b: out <= 1'b1;
24'h03802b: out <= 1'b1;
24'h03f02b: out <= 1'b1;
24'h04002b: out <= 1'b1;
24'h04102b: out <= 1'b1;
24'h04202b: out <= 1'b1;
24'h04302b: out <= 1'b1;
24'h04402b: out <= 1'b1;
24'h04502b: out <= 1'b1;
24'h04702b: out <= 1'b1;
24'h04802b: out <= 1'b1;
24'h04902b: out <= 1'b1;
24'h04a02b: out <= 1'b1;
24'h04b02b: out <= 1'b1;
24'h04c02b: out <= 1'b1;
24'h04d02b: out <= 1'b1;
24'h04e02b: out <= 1'b1;
24'h04f02b: out <= 1'b1;
24'h05002b: out <= 1'b1;
24'h05102b: out <= 1'b1;
24'h05202b: out <= 1'b1;
24'h05302b: out <= 1'b1;
24'h05402b: out <= 1'b1;
24'h05502b: out <= 1'b1;
24'h05602b: out <= 1'b1;
24'h05702b: out <= 1'b1;
24'h05802b: out <= 1'b1;
24'h05902b: out <= 1'b1;
24'h05a02b: out <= 1'b1;
24'h05b02b: out <= 1'b1;
24'h00b02c: out <= 1'b1;
24'h00c02c: out <= 1'b1;
24'h00d02c: out <= 1'b1;
24'h00e02c: out <= 1'b1;
24'h00f02c: out <= 1'b1;
24'h01002c: out <= 1'b1;
24'h01102c: out <= 1'b1;
24'h01202c: out <= 1'b1;
24'h01302c: out <= 1'b1;
24'h01402c: out <= 1'b1;
24'h01502c: out <= 1'b1;
24'h01602c: out <= 1'b1;
24'h01702c: out <= 1'b1;
24'h01802c: out <= 1'b1;
24'h01902c: out <= 1'b1;
24'h01c02c: out <= 1'b1;
24'h01d02c: out <= 1'b1;
24'h01e02c: out <= 1'b1;
24'h01f02c: out <= 1'b1;
24'h02002c: out <= 1'b1;
24'h02102c: out <= 1'b1;
24'h02202c: out <= 1'b1;
24'h02902c: out <= 1'b1;
24'h02a02c: out <= 1'b1;
24'h02b02c: out <= 1'b1;
24'h02c02c: out <= 1'b1;
24'h02d02c: out <= 1'b1;
24'h02e02c: out <= 1'b1;
24'h02f02c: out <= 1'b1;
24'h03202c: out <= 1'b1;
24'h03302c: out <= 1'b1;
24'h03402c: out <= 1'b1;
24'h03502c: out <= 1'b1;
24'h03602c: out <= 1'b1;
24'h03702c: out <= 1'b1;
24'h03802c: out <= 1'b1;
24'h03f02c: out <= 1'b1;
24'h04002c: out <= 1'b1;
24'h04102c: out <= 1'b1;
24'h04202c: out <= 1'b1;
24'h04302c: out <= 1'b1;
24'h04402c: out <= 1'b1;
24'h04502c: out <= 1'b1;
24'h04702c: out <= 1'b1;
24'h04802c: out <= 1'b1;
24'h04902c: out <= 1'b1;
24'h04a02c: out <= 1'b1;
24'h04b02c: out <= 1'b1;
24'h04c02c: out <= 1'b1;
24'h04d02c: out <= 1'b1;
24'h04e02c: out <= 1'b1;
24'h04f02c: out <= 1'b1;
24'h05002c: out <= 1'b1;
24'h05102c: out <= 1'b1;
24'h05202c: out <= 1'b1;
24'h05302c: out <= 1'b1;
24'h05402c: out <= 1'b1;
24'h05502c: out <= 1'b1;
24'h05602c: out <= 1'b1;
24'h05702c: out <= 1'b1;
24'h05802c: out <= 1'b1;
24'h05902c: out <= 1'b1;
24'h05a02c: out <= 1'b1;
24'h05b02c: out <= 1'b1;
24'h00b02d: out <= 1'b1;
24'h00c02d: out <= 1'b1;
24'h00d02d: out <= 1'b1;
24'h00e02d: out <= 1'b1;
24'h00f02d: out <= 1'b1;
24'h01002d: out <= 1'b1;
24'h01102d: out <= 1'b1;
24'h01202d: out <= 1'b1;
24'h01302d: out <= 1'b1;
24'h01402d: out <= 1'b1;
24'h01502d: out <= 1'b1;
24'h01602d: out <= 1'b1;
24'h01702d: out <= 1'b1;
24'h01802d: out <= 1'b1;
24'h01902d: out <= 1'b1;
24'h01c02d: out <= 1'b1;
24'h01d02d: out <= 1'b1;
24'h01e02d: out <= 1'b1;
24'h01f02d: out <= 1'b1;
24'h02002d: out <= 1'b1;
24'h02102d: out <= 1'b1;
24'h02202d: out <= 1'b1;
24'h02902d: out <= 1'b1;
24'h02a02d: out <= 1'b1;
24'h02b02d: out <= 1'b1;
24'h02c02d: out <= 1'b1;
24'h02d02d: out <= 1'b1;
24'h02e02d: out <= 1'b1;
24'h02f02d: out <= 1'b1;
24'h03202d: out <= 1'b1;
24'h03302d: out <= 1'b1;
24'h03402d: out <= 1'b1;
24'h03502d: out <= 1'b1;
24'h03602d: out <= 1'b1;
24'h03702d: out <= 1'b1;
24'h03802d: out <= 1'b1;
24'h03f02d: out <= 1'b1;
24'h04002d: out <= 1'b1;
24'h04102d: out <= 1'b1;
24'h04202d: out <= 1'b1;
24'h04302d: out <= 1'b1;
24'h04402d: out <= 1'b1;
24'h04502d: out <= 1'b1;
24'h04702d: out <= 1'b1;
24'h04802d: out <= 1'b1;
24'h04902d: out <= 1'b1;
24'h04a02d: out <= 1'b1;
24'h04b02d: out <= 1'b1;
24'h04c02d: out <= 1'b1;
24'h04d02d: out <= 1'b1;
24'h04e02d: out <= 1'b1;
24'h04f02d: out <= 1'b1;
24'h05002d: out <= 1'b1;
24'h05102d: out <= 1'b1;
24'h05202d: out <= 1'b1;
24'h05302d: out <= 1'b1;
24'h05402d: out <= 1'b1;
24'h05502d: out <= 1'b1;
24'h05602d: out <= 1'b1;
24'h05702d: out <= 1'b1;
24'h05802d: out <= 1'b1;
24'h05902d: out <= 1'b1;
24'h05a02d: out <= 1'b1;
24'h05b02d: out <= 1'b1;
24'h00c02e: out <= 1'b1;
24'h00d02e: out <= 1'b1;
24'h00e02e: out <= 1'b1;
24'h00f02e: out <= 1'b1;
24'h01002e: out <= 1'b1;
24'h01102e: out <= 1'b1;
24'h01202e: out <= 1'b1;
24'h01302e: out <= 1'b1;
24'h01402e: out <= 1'b1;
24'h01502e: out <= 1'b1;
24'h01602e: out <= 1'b1;
24'h01702e: out <= 1'b1;
24'h01802e: out <= 1'b1;
24'h01902e: out <= 1'b1;
24'h01c02e: out <= 1'b1;
24'h01d02e: out <= 1'b1;
24'h01e02e: out <= 1'b1;
24'h01f02e: out <= 1'b1;
24'h02002e: out <= 1'b1;
24'h02102e: out <= 1'b1;
24'h02a02e: out <= 1'b1;
24'h02b02e: out <= 1'b1;
24'h02c02e: out <= 1'b1;
24'h02d02e: out <= 1'b1;
24'h02e02e: out <= 1'b1;
24'h03202e: out <= 1'b1;
24'h03302e: out <= 1'b1;
24'h03402e: out <= 1'b1;
24'h03502e: out <= 1'b1;
24'h03602e: out <= 1'b1;
24'h03702e: out <= 1'b1;
24'h03f02e: out <= 1'b1;
24'h04002e: out <= 1'b1;
24'h04102e: out <= 1'b1;
24'h04202e: out <= 1'b1;
24'h04302e: out <= 1'b1;
24'h04402e: out <= 1'b1;
24'h04802e: out <= 1'b1;
24'h04902e: out <= 1'b1;
24'h04a02e: out <= 1'b1;
24'h04b02e: out <= 1'b1;
24'h04c02e: out <= 1'b1;
24'h04d02e: out <= 1'b1;
24'h04e02e: out <= 1'b1;
24'h04f02e: out <= 1'b1;
24'h05002e: out <= 1'b1;
24'h05102e: out <= 1'b1;
24'h05202e: out <= 1'b1;
24'h05302e: out <= 1'b1;
24'h05402e: out <= 1'b1;
24'h05502e: out <= 1'b1;
24'h05602e: out <= 1'b1;
24'h05702e: out <= 1'b1;
24'h05802e: out <= 1'b1;
24'h05902e: out <= 1'b1;
24'h05a02e: out <= 1'b1;
24'h009034: out <= 1'b1;
24'h00a034: out <= 1'b1;
24'h00b034: out <= 1'b1;
24'h00c034: out <= 1'b1;
24'h00d034: out <= 1'b1;
24'h00e034: out <= 1'b1;
24'h00f034: out <= 1'b1;
24'h010034: out <= 1'b1;
24'h011034: out <= 1'b1;
24'h012034: out <= 1'b1;
24'h013034: out <= 1'b1;
24'h014034: out <= 1'b1;
24'h015034: out <= 1'b1;
24'h016034: out <= 1'b1;
24'h01c034: out <= 1'b1;
24'h01d034: out <= 1'b1;
24'h01e034: out <= 1'b1;
24'h01f034: out <= 1'b1;
24'h020034: out <= 1'b1;
24'h021034: out <= 1'b1;
24'h022034: out <= 1'b1;
24'h029034: out <= 1'b1;
24'h02a034: out <= 1'b1;
24'h02b034: out <= 1'b1;
24'h02c034: out <= 1'b1;
24'h02d034: out <= 1'b1;
24'h02e034: out <= 1'b1;
24'h02f034: out <= 1'b1;
24'h032034: out <= 1'b1;
24'h033034: out <= 1'b1;
24'h034034: out <= 1'b1;
24'h035034: out <= 1'b1;
24'h036034: out <= 1'b1;
24'h037034: out <= 1'b1;
24'h038034: out <= 1'b1;
24'h039034: out <= 1'b1;
24'h03a034: out <= 1'b1;
24'h03b034: out <= 1'b1;
24'h03c034: out <= 1'b1;
24'h03d034: out <= 1'b1;
24'h03e034: out <= 1'b1;
24'h03f034: out <= 1'b1;
24'h040034: out <= 1'b1;
24'h041034: out <= 1'b1;
24'h042034: out <= 1'b1;
24'h043034: out <= 1'b1;
24'h044034: out <= 1'b1;
24'h045034: out <= 1'b1;
24'h048034: out <= 1'b1;
24'h049034: out <= 1'b1;
24'h04a034: out <= 1'b1;
24'h04b034: out <= 1'b1;
24'h04c034: out <= 1'b1;
24'h04d034: out <= 1'b1;
24'h04e034: out <= 1'b1;
24'h04f034: out <= 1'b1;
24'h050034: out <= 1'b1;
24'h051034: out <= 1'b1;
24'h052034: out <= 1'b1;
24'h053034: out <= 1'b1;
24'h054034: out <= 1'b1;
24'h055034: out <= 1'b1;
24'h056034: out <= 1'b1;
24'h057034: out <= 1'b1;
24'h058034: out <= 1'b1;
24'h008035: out <= 1'b1;
24'h009035: out <= 1'b1;
24'h00a035: out <= 1'b1;
24'h00b035: out <= 1'b1;
24'h00c035: out <= 1'b1;
24'h00d035: out <= 1'b1;
24'h00e035: out <= 1'b1;
24'h00f035: out <= 1'b1;
24'h010035: out <= 1'b1;
24'h011035: out <= 1'b1;
24'h012035: out <= 1'b1;
24'h013035: out <= 1'b1;
24'h014035: out <= 1'b1;
24'h015035: out <= 1'b1;
24'h016035: out <= 1'b1;
24'h01c035: out <= 1'b1;
24'h01d035: out <= 1'b1;
24'h01e035: out <= 1'b1;
24'h01f035: out <= 1'b1;
24'h020035: out <= 1'b1;
24'h021035: out <= 1'b1;
24'h022035: out <= 1'b1;
24'h029035: out <= 1'b1;
24'h02a035: out <= 1'b1;
24'h02b035: out <= 1'b1;
24'h02c035: out <= 1'b1;
24'h02d035: out <= 1'b1;
24'h02e035: out <= 1'b1;
24'h02f035: out <= 1'b1;
24'h032035: out <= 1'b1;
24'h033035: out <= 1'b1;
24'h034035: out <= 1'b1;
24'h035035: out <= 1'b1;
24'h036035: out <= 1'b1;
24'h037035: out <= 1'b1;
24'h038035: out <= 1'b1;
24'h039035: out <= 1'b1;
24'h03a035: out <= 1'b1;
24'h03b035: out <= 1'b1;
24'h03c035: out <= 1'b1;
24'h03d035: out <= 1'b1;
24'h03e035: out <= 1'b1;
24'h03f035: out <= 1'b1;
24'h040035: out <= 1'b1;
24'h041035: out <= 1'b1;
24'h042035: out <= 1'b1;
24'h043035: out <= 1'b1;
24'h044035: out <= 1'b1;
24'h045035: out <= 1'b1;
24'h047035: out <= 1'b1;
24'h048035: out <= 1'b1;
24'h049035: out <= 1'b1;
24'h04a035: out <= 1'b1;
24'h04b035: out <= 1'b1;
24'h04c035: out <= 1'b1;
24'h04d035: out <= 1'b1;
24'h04e035: out <= 1'b1;
24'h04f035: out <= 1'b1;
24'h050035: out <= 1'b1;
24'h051035: out <= 1'b1;
24'h052035: out <= 1'b1;
24'h053035: out <= 1'b1;
24'h054035: out <= 1'b1;
24'h055035: out <= 1'b1;
24'h056035: out <= 1'b1;
24'h057035: out <= 1'b1;
24'h058035: out <= 1'b1;
24'h007036: out <= 1'b1;
24'h008036: out <= 1'b1;
24'h009036: out <= 1'b1;
24'h00a036: out <= 1'b1;
24'h00b036: out <= 1'b1;
24'h00c036: out <= 1'b1;
24'h00d036: out <= 1'b1;
24'h00e036: out <= 1'b1;
24'h00f036: out <= 1'b1;
24'h010036: out <= 1'b1;
24'h011036: out <= 1'b1;
24'h012036: out <= 1'b1;
24'h013036: out <= 1'b1;
24'h014036: out <= 1'b1;
24'h015036: out <= 1'b1;
24'h016036: out <= 1'b1;
24'h017036: out <= 1'b1;
24'h018036: out <= 1'b1;
24'h01c036: out <= 1'b1;
24'h01d036: out <= 1'b1;
24'h01e036: out <= 1'b1;
24'h01f036: out <= 1'b1;
24'h020036: out <= 1'b1;
24'h021036: out <= 1'b1;
24'h022036: out <= 1'b1;
24'h029036: out <= 1'b1;
24'h02a036: out <= 1'b1;
24'h02b036: out <= 1'b1;
24'h02c036: out <= 1'b1;
24'h02d036: out <= 1'b1;
24'h02e036: out <= 1'b1;
24'h02f036: out <= 1'b1;
24'h032036: out <= 1'b1;
24'h033036: out <= 1'b1;
24'h034036: out <= 1'b1;
24'h035036: out <= 1'b1;
24'h036036: out <= 1'b1;
24'h037036: out <= 1'b1;
24'h038036: out <= 1'b1;
24'h039036: out <= 1'b1;
24'h03a036: out <= 1'b1;
24'h03b036: out <= 1'b1;
24'h03c036: out <= 1'b1;
24'h03d036: out <= 1'b1;
24'h03e036: out <= 1'b1;
24'h03f036: out <= 1'b1;
24'h040036: out <= 1'b1;
24'h041036: out <= 1'b1;
24'h042036: out <= 1'b1;
24'h043036: out <= 1'b1;
24'h044036: out <= 1'b1;
24'h045036: out <= 1'b1;
24'h047036: out <= 1'b1;
24'h048036: out <= 1'b1;
24'h049036: out <= 1'b1;
24'h04a036: out <= 1'b1;
24'h04b036: out <= 1'b1;
24'h04c036: out <= 1'b1;
24'h04d036: out <= 1'b1;
24'h04e036: out <= 1'b1;
24'h04f036: out <= 1'b1;
24'h050036: out <= 1'b1;
24'h051036: out <= 1'b1;
24'h052036: out <= 1'b1;
24'h053036: out <= 1'b1;
24'h054036: out <= 1'b1;
24'h055036: out <= 1'b1;
24'h056036: out <= 1'b1;
24'h057036: out <= 1'b1;
24'h058036: out <= 1'b1;
24'h059036: out <= 1'b1;
24'h05a036: out <= 1'b1;
24'h006037: out <= 1'b1;
24'h007037: out <= 1'b1;
24'h008037: out <= 1'b1;
24'h009037: out <= 1'b1;
24'h00a037: out <= 1'b1;
24'h00b037: out <= 1'b1;
24'h00c037: out <= 1'b1;
24'h00d037: out <= 1'b1;
24'h00e037: out <= 1'b1;
24'h00f037: out <= 1'b1;
24'h010037: out <= 1'b1;
24'h011037: out <= 1'b1;
24'h012037: out <= 1'b1;
24'h013037: out <= 1'b1;
24'h014037: out <= 1'b1;
24'h015037: out <= 1'b1;
24'h016037: out <= 1'b1;
24'h017037: out <= 1'b1;
24'h018037: out <= 1'b1;
24'h019037: out <= 1'b1;
24'h01c037: out <= 1'b1;
24'h01d037: out <= 1'b1;
24'h01e037: out <= 1'b1;
24'h01f037: out <= 1'b1;
24'h020037: out <= 1'b1;
24'h021037: out <= 1'b1;
24'h022037: out <= 1'b1;
24'h029037: out <= 1'b1;
24'h02a037: out <= 1'b1;
24'h02b037: out <= 1'b1;
24'h02c037: out <= 1'b1;
24'h02d037: out <= 1'b1;
24'h02e037: out <= 1'b1;
24'h02f037: out <= 1'b1;
24'h032037: out <= 1'b1;
24'h033037: out <= 1'b1;
24'h034037: out <= 1'b1;
24'h035037: out <= 1'b1;
24'h036037: out <= 1'b1;
24'h037037: out <= 1'b1;
24'h038037: out <= 1'b1;
24'h039037: out <= 1'b1;
24'h03a037: out <= 1'b1;
24'h03b037: out <= 1'b1;
24'h03c037: out <= 1'b1;
24'h03d037: out <= 1'b1;
24'h03e037: out <= 1'b1;
24'h03f037: out <= 1'b1;
24'h040037: out <= 1'b1;
24'h041037: out <= 1'b1;
24'h042037: out <= 1'b1;
24'h043037: out <= 1'b1;
24'h044037: out <= 1'b1;
24'h045037: out <= 1'b1;
24'h047037: out <= 1'b1;
24'h048037: out <= 1'b1;
24'h049037: out <= 1'b1;
24'h04a037: out <= 1'b1;
24'h04b037: out <= 1'b1;
24'h04c037: out <= 1'b1;
24'h04d037: out <= 1'b1;
24'h04e037: out <= 1'b1;
24'h04f037: out <= 1'b1;
24'h050037: out <= 1'b1;
24'h051037: out <= 1'b1;
24'h052037: out <= 1'b1;
24'h053037: out <= 1'b1;
24'h054037: out <= 1'b1;
24'h055037: out <= 1'b1;
24'h056037: out <= 1'b1;
24'h057037: out <= 1'b1;
24'h058037: out <= 1'b1;
24'h059037: out <= 1'b1;
24'h05a037: out <= 1'b1;
24'h05b037: out <= 1'b1;
24'h006038: out <= 1'b1;
24'h007038: out <= 1'b1;
24'h008038: out <= 1'b1;
24'h009038: out <= 1'b1;
24'h00a038: out <= 1'b1;
24'h00b038: out <= 1'b1;
24'h00c038: out <= 1'b1;
24'h013038: out <= 1'b1;
24'h014038: out <= 1'b1;
24'h015038: out <= 1'b1;
24'h016038: out <= 1'b1;
24'h017038: out <= 1'b1;
24'h018038: out <= 1'b1;
24'h019038: out <= 1'b1;
24'h01c038: out <= 1'b1;
24'h01d038: out <= 1'b1;
24'h01e038: out <= 1'b1;
24'h01f038: out <= 1'b1;
24'h020038: out <= 1'b1;
24'h021038: out <= 1'b1;
24'h022038: out <= 1'b1;
24'h029038: out <= 1'b1;
24'h02a038: out <= 1'b1;
24'h02b038: out <= 1'b1;
24'h02c038: out <= 1'b1;
24'h02d038: out <= 1'b1;
24'h02e038: out <= 1'b1;
24'h02f038: out <= 1'b1;
24'h032038: out <= 1'b1;
24'h033038: out <= 1'b1;
24'h034038: out <= 1'b1;
24'h035038: out <= 1'b1;
24'h036038: out <= 1'b1;
24'h037038: out <= 1'b1;
24'h038038: out <= 1'b1;
24'h047038: out <= 1'b1;
24'h048038: out <= 1'b1;
24'h049038: out <= 1'b1;
24'h04a038: out <= 1'b1;
24'h04b038: out <= 1'b1;
24'h04c038: out <= 1'b1;
24'h04d038: out <= 1'b1;
24'h04e038: out <= 1'b1;
24'h055038: out <= 1'b1;
24'h056038: out <= 1'b1;
24'h057038: out <= 1'b1;
24'h058038: out <= 1'b1;
24'h059038: out <= 1'b1;
24'h05a038: out <= 1'b1;
24'h05b038: out <= 1'b1;
24'h006039: out <= 1'b1;
24'h007039: out <= 1'b1;
24'h008039: out <= 1'b1;
24'h009039: out <= 1'b1;
24'h00a039: out <= 1'b1;
24'h00b039: out <= 1'b1;
24'h00c039: out <= 1'b1;
24'h013039: out <= 1'b1;
24'h014039: out <= 1'b1;
24'h015039: out <= 1'b1;
24'h016039: out <= 1'b1;
24'h017039: out <= 1'b1;
24'h018039: out <= 1'b1;
24'h019039: out <= 1'b1;
24'h01c039: out <= 1'b1;
24'h01d039: out <= 1'b1;
24'h01e039: out <= 1'b1;
24'h01f039: out <= 1'b1;
24'h020039: out <= 1'b1;
24'h021039: out <= 1'b1;
24'h022039: out <= 1'b1;
24'h029039: out <= 1'b1;
24'h02a039: out <= 1'b1;
24'h02b039: out <= 1'b1;
24'h02c039: out <= 1'b1;
24'h02d039: out <= 1'b1;
24'h02e039: out <= 1'b1;
24'h02f039: out <= 1'b1;
24'h032039: out <= 1'b1;
24'h033039: out <= 1'b1;
24'h034039: out <= 1'b1;
24'h035039: out <= 1'b1;
24'h036039: out <= 1'b1;
24'h037039: out <= 1'b1;
24'h038039: out <= 1'b1;
24'h047039: out <= 1'b1;
24'h048039: out <= 1'b1;
24'h049039: out <= 1'b1;
24'h04a039: out <= 1'b1;
24'h04b039: out <= 1'b1;
24'h04c039: out <= 1'b1;
24'h04d039: out <= 1'b1;
24'h04e039: out <= 1'b1;
24'h055039: out <= 1'b1;
24'h056039: out <= 1'b1;
24'h057039: out <= 1'b1;
24'h058039: out <= 1'b1;
24'h059039: out <= 1'b1;
24'h05a039: out <= 1'b1;
24'h05b039: out <= 1'b1;
24'h00603a: out <= 1'b1;
24'h00703a: out <= 1'b1;
24'h00803a: out <= 1'b1;
24'h00903a: out <= 1'b1;
24'h00a03a: out <= 1'b1;
24'h00b03a: out <= 1'b1;
24'h00c03a: out <= 1'b1;
24'h01303a: out <= 1'b1;
24'h01403a: out <= 1'b1;
24'h01503a: out <= 1'b1;
24'h01603a: out <= 1'b1;
24'h01703a: out <= 1'b1;
24'h01803a: out <= 1'b1;
24'h01903a: out <= 1'b1;
24'h01c03a: out <= 1'b1;
24'h01d03a: out <= 1'b1;
24'h01e03a: out <= 1'b1;
24'h01f03a: out <= 1'b1;
24'h02003a: out <= 1'b1;
24'h02103a: out <= 1'b1;
24'h02203a: out <= 1'b1;
24'h02903a: out <= 1'b1;
24'h02a03a: out <= 1'b1;
24'h02b03a: out <= 1'b1;
24'h02c03a: out <= 1'b1;
24'h02d03a: out <= 1'b1;
24'h02e03a: out <= 1'b1;
24'h02f03a: out <= 1'b1;
24'h03203a: out <= 1'b1;
24'h03303a: out <= 1'b1;
24'h03403a: out <= 1'b1;
24'h03503a: out <= 1'b1;
24'h03603a: out <= 1'b1;
24'h03703a: out <= 1'b1;
24'h03803a: out <= 1'b1;
24'h04703a: out <= 1'b1;
24'h04803a: out <= 1'b1;
24'h04903a: out <= 1'b1;
24'h04a03a: out <= 1'b1;
24'h04b03a: out <= 1'b1;
24'h04c03a: out <= 1'b1;
24'h04d03a: out <= 1'b1;
24'h04e03a: out <= 1'b1;
24'h05503a: out <= 1'b1;
24'h05603a: out <= 1'b1;
24'h05703a: out <= 1'b1;
24'h05803a: out <= 1'b1;
24'h05903a: out <= 1'b1;
24'h05a03a: out <= 1'b1;
24'h05b03a: out <= 1'b1;
24'h00603b: out <= 1'b1;
24'h00703b: out <= 1'b1;
24'h00803b: out <= 1'b1;
24'h00903b: out <= 1'b1;
24'h00a03b: out <= 1'b1;
24'h00b03b: out <= 1'b1;
24'h00c03b: out <= 1'b1;
24'h01303b: out <= 1'b1;
24'h01403b: out <= 1'b1;
24'h01503b: out <= 1'b1;
24'h01603b: out <= 1'b1;
24'h01703b: out <= 1'b1;
24'h01803b: out <= 1'b1;
24'h01903b: out <= 1'b1;
24'h01c03b: out <= 1'b1;
24'h01d03b: out <= 1'b1;
24'h01e03b: out <= 1'b1;
24'h01f03b: out <= 1'b1;
24'h02003b: out <= 1'b1;
24'h02103b: out <= 1'b1;
24'h02203b: out <= 1'b1;
24'h02903b: out <= 1'b1;
24'h02a03b: out <= 1'b1;
24'h02b03b: out <= 1'b1;
24'h02c03b: out <= 1'b1;
24'h02d03b: out <= 1'b1;
24'h02e03b: out <= 1'b1;
24'h02f03b: out <= 1'b1;
24'h03203b: out <= 1'b1;
24'h03303b: out <= 1'b1;
24'h03403b: out <= 1'b1;
24'h03503b: out <= 1'b1;
24'h03603b: out <= 1'b1;
24'h03703b: out <= 1'b1;
24'h03803b: out <= 1'b1;
24'h04703b: out <= 1'b1;
24'h04803b: out <= 1'b1;
24'h04903b: out <= 1'b1;
24'h04a03b: out <= 1'b1;
24'h04b03b: out <= 1'b1;
24'h04c03b: out <= 1'b1;
24'h04d03b: out <= 1'b1;
24'h04e03b: out <= 1'b1;
24'h05503b: out <= 1'b1;
24'h05603b: out <= 1'b1;
24'h05703b: out <= 1'b1;
24'h05803b: out <= 1'b1;
24'h05903b: out <= 1'b1;
24'h05a03b: out <= 1'b1;
24'h05b03b: out <= 1'b1;
24'h00603c: out <= 1'b1;
24'h00703c: out <= 1'b1;
24'h00803c: out <= 1'b1;
24'h00903c: out <= 1'b1;
24'h00a03c: out <= 1'b1;
24'h00b03c: out <= 1'b1;
24'h00c03c: out <= 1'b1;
24'h01303c: out <= 1'b1;
24'h01403c: out <= 1'b1;
24'h01503c: out <= 1'b1;
24'h01603c: out <= 1'b1;
24'h01703c: out <= 1'b1;
24'h01803c: out <= 1'b1;
24'h01903c: out <= 1'b1;
24'h01c03c: out <= 1'b1;
24'h01d03c: out <= 1'b1;
24'h01e03c: out <= 1'b1;
24'h01f03c: out <= 1'b1;
24'h02003c: out <= 1'b1;
24'h02103c: out <= 1'b1;
24'h02203c: out <= 1'b1;
24'h02303c: out <= 1'b1;
24'h02403c: out <= 1'b1;
24'h02603c: out <= 1'b1;
24'h02703c: out <= 1'b1;
24'h02803c: out <= 1'b1;
24'h02903c: out <= 1'b1;
24'h02a03c: out <= 1'b1;
24'h02b03c: out <= 1'b1;
24'h02c03c: out <= 1'b1;
24'h02d03c: out <= 1'b1;
24'h02e03c: out <= 1'b1;
24'h02f03c: out <= 1'b1;
24'h03203c: out <= 1'b1;
24'h03303c: out <= 1'b1;
24'h03403c: out <= 1'b1;
24'h03503c: out <= 1'b1;
24'h03603c: out <= 1'b1;
24'h03703c: out <= 1'b1;
24'h03803c: out <= 1'b1;
24'h03903c: out <= 1'b1;
24'h03a03c: out <= 1'b1;
24'h03b03c: out <= 1'b1;
24'h03c03c: out <= 1'b1;
24'h03d03c: out <= 1'b1;
24'h03e03c: out <= 1'b1;
24'h03f03c: out <= 1'b1;
24'h04003c: out <= 1'b1;
24'h04103c: out <= 1'b1;
24'h04203c: out <= 1'b1;
24'h04703c: out <= 1'b1;
24'h04803c: out <= 1'b1;
24'h04903c: out <= 1'b1;
24'h04a03c: out <= 1'b1;
24'h04b03c: out <= 1'b1;
24'h04c03c: out <= 1'b1;
24'h04d03c: out <= 1'b1;
24'h04e03c: out <= 1'b1;
24'h05203c: out <= 1'b1;
24'h05303c: out <= 1'b1;
24'h05403c: out <= 1'b1;
24'h05503c: out <= 1'b1;
24'h05603c: out <= 1'b1;
24'h05703c: out <= 1'b1;
24'h05803c: out <= 1'b1;
24'h05903c: out <= 1'b1;
24'h05a03c: out <= 1'b1;
24'h05b03c: out <= 1'b1;
24'h00603d: out <= 1'b1;
24'h00703d: out <= 1'b1;
24'h00803d: out <= 1'b1;
24'h00903d: out <= 1'b1;
24'h00a03d: out <= 1'b1;
24'h00b03d: out <= 1'b1;
24'h00c03d: out <= 1'b1;
24'h01303d: out <= 1'b1;
24'h01403d: out <= 1'b1;
24'h01503d: out <= 1'b1;
24'h01603d: out <= 1'b1;
24'h01703d: out <= 1'b1;
24'h01803d: out <= 1'b1;
24'h01903d: out <= 1'b1;
24'h01c03d: out <= 1'b1;
24'h01d03d: out <= 1'b1;
24'h01e03d: out <= 1'b1;
24'h01f03d: out <= 1'b1;
24'h02003d: out <= 1'b1;
24'h02103d: out <= 1'b1;
24'h02203d: out <= 1'b1;
24'h02303d: out <= 1'b1;
24'h02403d: out <= 1'b1;
24'h02603d: out <= 1'b1;
24'h02703d: out <= 1'b1;
24'h02803d: out <= 1'b1;
24'h02903d: out <= 1'b1;
24'h02a03d: out <= 1'b1;
24'h02b03d: out <= 1'b1;
24'h02c03d: out <= 1'b1;
24'h02d03d: out <= 1'b1;
24'h02e03d: out <= 1'b1;
24'h02f03d: out <= 1'b1;
24'h03203d: out <= 1'b1;
24'h03303d: out <= 1'b1;
24'h03403d: out <= 1'b1;
24'h03503d: out <= 1'b1;
24'h03603d: out <= 1'b1;
24'h03703d: out <= 1'b1;
24'h03803d: out <= 1'b1;
24'h03903d: out <= 1'b1;
24'h03a03d: out <= 1'b1;
24'h03b03d: out <= 1'b1;
24'h03c03d: out <= 1'b1;
24'h03d03d: out <= 1'b1;
24'h03e03d: out <= 1'b1;
24'h03f03d: out <= 1'b1;
24'h04003d: out <= 1'b1;
24'h04103d: out <= 1'b1;
24'h04203d: out <= 1'b1;
24'h04703d: out <= 1'b1;
24'h04803d: out <= 1'b1;
24'h04903d: out <= 1'b1;
24'h04a03d: out <= 1'b1;
24'h04b03d: out <= 1'b1;
24'h04c03d: out <= 1'b1;
24'h04d03d: out <= 1'b1;
24'h04e03d: out <= 1'b1;
24'h05203d: out <= 1'b1;
24'h05303d: out <= 1'b1;
24'h05403d: out <= 1'b1;
24'h05503d: out <= 1'b1;
24'h05603d: out <= 1'b1;
24'h05703d: out <= 1'b1;
24'h05803d: out <= 1'b1;
24'h05903d: out <= 1'b1;
24'h05a03d: out <= 1'b1;
24'h05b03d: out <= 1'b1;
24'h00603e: out <= 1'b1;
24'h00703e: out <= 1'b1;
24'h00803e: out <= 1'b1;
24'h00903e: out <= 1'b1;
24'h00a03e: out <= 1'b1;
24'h00b03e: out <= 1'b1;
24'h00c03e: out <= 1'b1;
24'h01303e: out <= 1'b1;
24'h01403e: out <= 1'b1;
24'h01503e: out <= 1'b1;
24'h01603e: out <= 1'b1;
24'h01703e: out <= 1'b1;
24'h01803e: out <= 1'b1;
24'h01903e: out <= 1'b1;
24'h01c03e: out <= 1'b1;
24'h01d03e: out <= 1'b1;
24'h01e03e: out <= 1'b1;
24'h01f03e: out <= 1'b1;
24'h02003e: out <= 1'b1;
24'h02103e: out <= 1'b1;
24'h02203e: out <= 1'b1;
24'h02303e: out <= 1'b1;
24'h02403e: out <= 1'b1;
24'h02503e: out <= 1'b1;
24'h02603e: out <= 1'b1;
24'h02703e: out <= 1'b1;
24'h02803e: out <= 1'b1;
24'h02903e: out <= 1'b1;
24'h02a03e: out <= 1'b1;
24'h02b03e: out <= 1'b1;
24'h02c03e: out <= 1'b1;
24'h02d03e: out <= 1'b1;
24'h02e03e: out <= 1'b1;
24'h02f03e: out <= 1'b1;
24'h03203e: out <= 1'b1;
24'h03303e: out <= 1'b1;
24'h03403e: out <= 1'b1;
24'h03503e: out <= 1'b1;
24'h03603e: out <= 1'b1;
24'h03703e: out <= 1'b1;
24'h03803e: out <= 1'b1;
24'h03903e: out <= 1'b1;
24'h03a03e: out <= 1'b1;
24'h03b03e: out <= 1'b1;
24'h03c03e: out <= 1'b1;
24'h03d03e: out <= 1'b1;
24'h03e03e: out <= 1'b1;
24'h03f03e: out <= 1'b1;
24'h04003e: out <= 1'b1;
24'h04103e: out <= 1'b1;
24'h04203e: out <= 1'b1;
24'h04703e: out <= 1'b1;
24'h04803e: out <= 1'b1;
24'h04903e: out <= 1'b1;
24'h04a03e: out <= 1'b1;
24'h04b03e: out <= 1'b1;
24'h04c03e: out <= 1'b1;
24'h04d03e: out <= 1'b1;
24'h04e03e: out <= 1'b1;
24'h04f03e: out <= 1'b1;
24'h05003e: out <= 1'b1;
24'h05103e: out <= 1'b1;
24'h05203e: out <= 1'b1;
24'h05303e: out <= 1'b1;
24'h05403e: out <= 1'b1;
24'h05503e: out <= 1'b1;
24'h05603e: out <= 1'b1;
24'h05703e: out <= 1'b1;
24'h05803e: out <= 1'b1;
24'h05903e: out <= 1'b1;
24'h05a03e: out <= 1'b1;
24'h05b03e: out <= 1'b1;
24'h00603f: out <= 1'b1;
24'h00703f: out <= 1'b1;
24'h00803f: out <= 1'b1;
24'h00903f: out <= 1'b1;
24'h00a03f: out <= 1'b1;
24'h00b03f: out <= 1'b1;
24'h00c03f: out <= 1'b1;
24'h01303f: out <= 1'b1;
24'h01403f: out <= 1'b1;
24'h01503f: out <= 1'b1;
24'h01603f: out <= 1'b1;
24'h01703f: out <= 1'b1;
24'h01803f: out <= 1'b1;
24'h01903f: out <= 1'b1;
24'h01c03f: out <= 1'b1;
24'h01d03f: out <= 1'b1;
24'h01e03f: out <= 1'b1;
24'h01f03f: out <= 1'b1;
24'h02003f: out <= 1'b1;
24'h02103f: out <= 1'b1;
24'h02203f: out <= 1'b1;
24'h02303f: out <= 1'b1;
24'h02403f: out <= 1'b1;
24'h02503f: out <= 1'b1;
24'h02603f: out <= 1'b1;
24'h02703f: out <= 1'b1;
24'h02803f: out <= 1'b1;
24'h02903f: out <= 1'b1;
24'h02a03f: out <= 1'b1;
24'h02b03f: out <= 1'b1;
24'h02c03f: out <= 1'b1;
24'h02d03f: out <= 1'b1;
24'h02e03f: out <= 1'b1;
24'h02f03f: out <= 1'b1;
24'h03203f: out <= 1'b1;
24'h03303f: out <= 1'b1;
24'h03403f: out <= 1'b1;
24'h03503f: out <= 1'b1;
24'h03603f: out <= 1'b1;
24'h03703f: out <= 1'b1;
24'h03803f: out <= 1'b1;
24'h03903f: out <= 1'b1;
24'h03a03f: out <= 1'b1;
24'h03b03f: out <= 1'b1;
24'h03c03f: out <= 1'b1;
24'h03d03f: out <= 1'b1;
24'h03e03f: out <= 1'b1;
24'h03f03f: out <= 1'b1;
24'h04003f: out <= 1'b1;
24'h04103f: out <= 1'b1;
24'h04203f: out <= 1'b1;
24'h04703f: out <= 1'b1;
24'h04803f: out <= 1'b1;
24'h04903f: out <= 1'b1;
24'h04a03f: out <= 1'b1;
24'h04b03f: out <= 1'b1;
24'h04c03f: out <= 1'b1;
24'h04d03f: out <= 1'b1;
24'h04e03f: out <= 1'b1;
24'h04f03f: out <= 1'b1;
24'h05003f: out <= 1'b1;
24'h05103f: out <= 1'b1;
24'h05203f: out <= 1'b1;
24'h05303f: out <= 1'b1;
24'h05403f: out <= 1'b1;
24'h05503f: out <= 1'b1;
24'h05603f: out <= 1'b1;
24'h05703f: out <= 1'b1;
24'h05803f: out <= 1'b1;
24'h05903f: out <= 1'b1;
24'h05a03f: out <= 1'b1;
24'h05b03f: out <= 1'b1;
24'h006040: out <= 1'b1;
24'h007040: out <= 1'b1;
24'h008040: out <= 1'b1;
24'h009040: out <= 1'b1;
24'h00a040: out <= 1'b1;
24'h00b040: out <= 1'b1;
24'h00c040: out <= 1'b1;
24'h013040: out <= 1'b1;
24'h014040: out <= 1'b1;
24'h015040: out <= 1'b1;
24'h016040: out <= 1'b1;
24'h017040: out <= 1'b1;
24'h018040: out <= 1'b1;
24'h019040: out <= 1'b1;
24'h01e040: out <= 1'b1;
24'h01f040: out <= 1'b1;
24'h020040: out <= 1'b1;
24'h021040: out <= 1'b1;
24'h022040: out <= 1'b1;
24'h023040: out <= 1'b1;
24'h024040: out <= 1'b1;
24'h025040: out <= 1'b1;
24'h026040: out <= 1'b1;
24'h027040: out <= 1'b1;
24'h028040: out <= 1'b1;
24'h029040: out <= 1'b1;
24'h02a040: out <= 1'b1;
24'h02b040: out <= 1'b1;
24'h02c040: out <= 1'b1;
24'h032040: out <= 1'b1;
24'h033040: out <= 1'b1;
24'h034040: out <= 1'b1;
24'h035040: out <= 1'b1;
24'h036040: out <= 1'b1;
24'h037040: out <= 1'b1;
24'h038040: out <= 1'b1;
24'h047040: out <= 1'b1;
24'h048040: out <= 1'b1;
24'h049040: out <= 1'b1;
24'h04a040: out <= 1'b1;
24'h04b040: out <= 1'b1;
24'h04c040: out <= 1'b1;
24'h04d040: out <= 1'b1;
24'h04e040: out <= 1'b1;
24'h04f040: out <= 1'b1;
24'h050040: out <= 1'b1;
24'h051040: out <= 1'b1;
24'h052040: out <= 1'b1;
24'h053040: out <= 1'b1;
24'h054040: out <= 1'b1;
24'h055040: out <= 1'b1;
24'h056040: out <= 1'b1;
24'h006041: out <= 1'b1;
24'h007041: out <= 1'b1;
24'h008041: out <= 1'b1;
24'h009041: out <= 1'b1;
24'h00a041: out <= 1'b1;
24'h00b041: out <= 1'b1;
24'h00c041: out <= 1'b1;
24'h013041: out <= 1'b1;
24'h014041: out <= 1'b1;
24'h015041: out <= 1'b1;
24'h016041: out <= 1'b1;
24'h017041: out <= 1'b1;
24'h018041: out <= 1'b1;
24'h019041: out <= 1'b1;
24'h01e041: out <= 1'b1;
24'h01f041: out <= 1'b1;
24'h020041: out <= 1'b1;
24'h021041: out <= 1'b1;
24'h022041: out <= 1'b1;
24'h023041: out <= 1'b1;
24'h024041: out <= 1'b1;
24'h025041: out <= 1'b1;
24'h026041: out <= 1'b1;
24'h027041: out <= 1'b1;
24'h028041: out <= 1'b1;
24'h029041: out <= 1'b1;
24'h02a041: out <= 1'b1;
24'h02b041: out <= 1'b1;
24'h02c041: out <= 1'b1;
24'h032041: out <= 1'b1;
24'h033041: out <= 1'b1;
24'h034041: out <= 1'b1;
24'h035041: out <= 1'b1;
24'h036041: out <= 1'b1;
24'h037041: out <= 1'b1;
24'h038041: out <= 1'b1;
24'h047041: out <= 1'b1;
24'h048041: out <= 1'b1;
24'h049041: out <= 1'b1;
24'h04a041: out <= 1'b1;
24'h04b041: out <= 1'b1;
24'h04c041: out <= 1'b1;
24'h04d041: out <= 1'b1;
24'h04e041: out <= 1'b1;
24'h04f041: out <= 1'b1;
24'h050041: out <= 1'b1;
24'h051041: out <= 1'b1;
24'h052041: out <= 1'b1;
24'h053041: out <= 1'b1;
24'h054041: out <= 1'b1;
24'h055041: out <= 1'b1;
24'h056041: out <= 1'b1;
24'h057041: out <= 1'b1;
24'h058041: out <= 1'b1;
24'h006042: out <= 1'b1;
24'h007042: out <= 1'b1;
24'h008042: out <= 1'b1;
24'h009042: out <= 1'b1;
24'h00a042: out <= 1'b1;
24'h00b042: out <= 1'b1;
24'h00c042: out <= 1'b1;
24'h013042: out <= 1'b1;
24'h014042: out <= 1'b1;
24'h015042: out <= 1'b1;
24'h016042: out <= 1'b1;
24'h017042: out <= 1'b1;
24'h018042: out <= 1'b1;
24'h019042: out <= 1'b1;
24'h01f042: out <= 1'b1;
24'h020042: out <= 1'b1;
24'h021042: out <= 1'b1;
24'h022042: out <= 1'b1;
24'h023042: out <= 1'b1;
24'h024042: out <= 1'b1;
24'h025042: out <= 1'b1;
24'h026042: out <= 1'b1;
24'h027042: out <= 1'b1;
24'h028042: out <= 1'b1;
24'h029042: out <= 1'b1;
24'h02a042: out <= 1'b1;
24'h02b042: out <= 1'b1;
24'h02c042: out <= 1'b1;
24'h032042: out <= 1'b1;
24'h033042: out <= 1'b1;
24'h034042: out <= 1'b1;
24'h035042: out <= 1'b1;
24'h036042: out <= 1'b1;
24'h037042: out <= 1'b1;
24'h038042: out <= 1'b1;
24'h047042: out <= 1'b1;
24'h048042: out <= 1'b1;
24'h049042: out <= 1'b1;
24'h04a042: out <= 1'b1;
24'h04b042: out <= 1'b1;
24'h04c042: out <= 1'b1;
24'h04d042: out <= 1'b1;
24'h04e042: out <= 1'b1;
24'h04f042: out <= 1'b1;
24'h050042: out <= 1'b1;
24'h051042: out <= 1'b1;
24'h052042: out <= 1'b1;
24'h053042: out <= 1'b1;
24'h054042: out <= 1'b1;
24'h055042: out <= 1'b1;
24'h056042: out <= 1'b1;
24'h057042: out <= 1'b1;
24'h058042: out <= 1'b1;
24'h006043: out <= 1'b1;
24'h007043: out <= 1'b1;
24'h008043: out <= 1'b1;
24'h009043: out <= 1'b1;
24'h00a043: out <= 1'b1;
24'h00b043: out <= 1'b1;
24'h00c043: out <= 1'b1;
24'h013043: out <= 1'b1;
24'h014043: out <= 1'b1;
24'h015043: out <= 1'b1;
24'h016043: out <= 1'b1;
24'h017043: out <= 1'b1;
24'h018043: out <= 1'b1;
24'h019043: out <= 1'b1;
24'h021043: out <= 1'b1;
24'h022043: out <= 1'b1;
24'h023043: out <= 1'b1;
24'h024043: out <= 1'b1;
24'h025043: out <= 1'b1;
24'h026043: out <= 1'b1;
24'h027043: out <= 1'b1;
24'h028043: out <= 1'b1;
24'h029043: out <= 1'b1;
24'h02a043: out <= 1'b1;
24'h032043: out <= 1'b1;
24'h033043: out <= 1'b1;
24'h034043: out <= 1'b1;
24'h035043: out <= 1'b1;
24'h036043: out <= 1'b1;
24'h037043: out <= 1'b1;
24'h038043: out <= 1'b1;
24'h047043: out <= 1'b1;
24'h048043: out <= 1'b1;
24'h049043: out <= 1'b1;
24'h04a043: out <= 1'b1;
24'h04b043: out <= 1'b1;
24'h04c043: out <= 1'b1;
24'h04d043: out <= 1'b1;
24'h04e043: out <= 1'b1;
24'h04f043: out <= 1'b1;
24'h050043: out <= 1'b1;
24'h051043: out <= 1'b1;
24'h052043: out <= 1'b1;
24'h053043: out <= 1'b1;
24'h054043: out <= 1'b1;
24'h055043: out <= 1'b1;
24'h056043: out <= 1'b1;
24'h057043: out <= 1'b1;
24'h058043: out <= 1'b1;
24'h006044: out <= 1'b1;
24'h007044: out <= 1'b1;
24'h008044: out <= 1'b1;
24'h009044: out <= 1'b1;
24'h00a044: out <= 1'b1;
24'h00b044: out <= 1'b1;
24'h00c044: out <= 1'b1;
24'h00d044: out <= 1'b1;
24'h00e044: out <= 1'b1;
24'h00f044: out <= 1'b1;
24'h010044: out <= 1'b1;
24'h011044: out <= 1'b1;
24'h012044: out <= 1'b1;
24'h013044: out <= 1'b1;
24'h014044: out <= 1'b1;
24'h015044: out <= 1'b1;
24'h016044: out <= 1'b1;
24'h017044: out <= 1'b1;
24'h018044: out <= 1'b1;
24'h019044: out <= 1'b1;
24'h021044: out <= 1'b1;
24'h022044: out <= 1'b1;
24'h023044: out <= 1'b1;
24'h024044: out <= 1'b1;
24'h025044: out <= 1'b1;
24'h026044: out <= 1'b1;
24'h027044: out <= 1'b1;
24'h028044: out <= 1'b1;
24'h029044: out <= 1'b1;
24'h02a044: out <= 1'b1;
24'h032044: out <= 1'b1;
24'h033044: out <= 1'b1;
24'h034044: out <= 1'b1;
24'h035044: out <= 1'b1;
24'h036044: out <= 1'b1;
24'h037044: out <= 1'b1;
24'h038044: out <= 1'b1;
24'h039044: out <= 1'b1;
24'h03a044: out <= 1'b1;
24'h03b044: out <= 1'b1;
24'h03c044: out <= 1'b1;
24'h03d044: out <= 1'b1;
24'h03e044: out <= 1'b1;
24'h03f044: out <= 1'b1;
24'h040044: out <= 1'b1;
24'h041044: out <= 1'b1;
24'h042044: out <= 1'b1;
24'h043044: out <= 1'b1;
24'h044044: out <= 1'b1;
24'h045044: out <= 1'b1;
24'h047044: out <= 1'b1;
24'h048044: out <= 1'b1;
24'h049044: out <= 1'b1;
24'h04a044: out <= 1'b1;
24'h04b044: out <= 1'b1;
24'h04c044: out <= 1'b1;
24'h04d044: out <= 1'b1;
24'h04e044: out <= 1'b1;
24'h04f044: out <= 1'b1;
24'h050044: out <= 1'b1;
24'h051044: out <= 1'b1;
24'h052044: out <= 1'b1;
24'h053044: out <= 1'b1;
24'h054044: out <= 1'b1;
24'h055044: out <= 1'b1;
24'h056044: out <= 1'b1;
24'h057044: out <= 1'b1;
24'h058044: out <= 1'b1;
24'h059044: out <= 1'b1;
24'h05a044: out <= 1'b1;
24'h05b044: out <= 1'b1;
24'h007045: out <= 1'b1;
24'h008045: out <= 1'b1;
24'h009045: out <= 1'b1;
24'h00a045: out <= 1'b1;
24'h00b045: out <= 1'b1;
24'h00c045: out <= 1'b1;
24'h00d045: out <= 1'b1;
24'h00e045: out <= 1'b1;
24'h00f045: out <= 1'b1;
24'h010045: out <= 1'b1;
24'h011045: out <= 1'b1;
24'h012045: out <= 1'b1;
24'h013045: out <= 1'b1;
24'h014045: out <= 1'b1;
24'h015045: out <= 1'b1;
24'h016045: out <= 1'b1;
24'h017045: out <= 1'b1;
24'h018045: out <= 1'b1;
24'h022045: out <= 1'b1;
24'h023045: out <= 1'b1;
24'h024045: out <= 1'b1;
24'h025045: out <= 1'b1;
24'h026045: out <= 1'b1;
24'h027045: out <= 1'b1;
24'h028045: out <= 1'b1;
24'h029045: out <= 1'b1;
24'h032045: out <= 1'b1;
24'h033045: out <= 1'b1;
24'h034045: out <= 1'b1;
24'h035045: out <= 1'b1;
24'h036045: out <= 1'b1;
24'h037045: out <= 1'b1;
24'h038045: out <= 1'b1;
24'h039045: out <= 1'b1;
24'h03a045: out <= 1'b1;
24'h03b045: out <= 1'b1;
24'h03c045: out <= 1'b1;
24'h03d045: out <= 1'b1;
24'h03e045: out <= 1'b1;
24'h03f045: out <= 1'b1;
24'h040045: out <= 1'b1;
24'h041045: out <= 1'b1;
24'h042045: out <= 1'b1;
24'h043045: out <= 1'b1;
24'h044045: out <= 1'b1;
24'h045045: out <= 1'b1;
24'h047045: out <= 1'b1;
24'h048045: out <= 1'b1;
24'h049045: out <= 1'b1;
24'h04a045: out <= 1'b1;
24'h04b045: out <= 1'b1;
24'h04c045: out <= 1'b1;
24'h04d045: out <= 1'b1;
24'h04e045: out <= 1'b1;
24'h050045: out <= 1'b1;
24'h051045: out <= 1'b1;
24'h052045: out <= 1'b1;
24'h053045: out <= 1'b1;
24'h054045: out <= 1'b1;
24'h055045: out <= 1'b1;
24'h056045: out <= 1'b1;
24'h057045: out <= 1'b1;
24'h058045: out <= 1'b1;
24'h059045: out <= 1'b1;
24'h05a045: out <= 1'b1;
24'h05b045: out <= 1'b1;
24'h008046: out <= 1'b1;
24'h009046: out <= 1'b1;
24'h00a046: out <= 1'b1;
24'h00b046: out <= 1'b1;
24'h00c046: out <= 1'b1;
24'h00d046: out <= 1'b1;
24'h00e046: out <= 1'b1;
24'h00f046: out <= 1'b1;
24'h010046: out <= 1'b1;
24'h011046: out <= 1'b1;
24'h012046: out <= 1'b1;
24'h013046: out <= 1'b1;
24'h014046: out <= 1'b1;
24'h015046: out <= 1'b1;
24'h016046: out <= 1'b1;
24'h024046: out <= 1'b1;
24'h025046: out <= 1'b1;
24'h026046: out <= 1'b1;
24'h027046: out <= 1'b1;
24'h032046: out <= 1'b1;
24'h033046: out <= 1'b1;
24'h034046: out <= 1'b1;
24'h035046: out <= 1'b1;
24'h036046: out <= 1'b1;
24'h037046: out <= 1'b1;
24'h038046: out <= 1'b1;
24'h039046: out <= 1'b1;
24'h03a046: out <= 1'b1;
24'h03b046: out <= 1'b1;
24'h03c046: out <= 1'b1;
24'h03d046: out <= 1'b1;
24'h03e046: out <= 1'b1;
24'h03f046: out <= 1'b1;
24'h040046: out <= 1'b1;
24'h041046: out <= 1'b1;
24'h042046: out <= 1'b1;
24'h043046: out <= 1'b1;
24'h044046: out <= 1'b1;
24'h045046: out <= 1'b1;
24'h047046: out <= 1'b1;
24'h048046: out <= 1'b1;
24'h049046: out <= 1'b1;
24'h04a046: out <= 1'b1;
24'h04b046: out <= 1'b1;
24'h04c046: out <= 1'b1;
24'h04d046: out <= 1'b1;
24'h04e046: out <= 1'b1;
24'h052046: out <= 1'b1;
24'h053046: out <= 1'b1;
24'h054046: out <= 1'b1;
24'h055046: out <= 1'b1;
24'h056046: out <= 1'b1;
24'h057046: out <= 1'b1;
24'h058046: out <= 1'b1;
24'h059046: out <= 1'b1;
24'h05a046: out <= 1'b1;
24'h05b046: out <= 1'b1;
24'h009047: out <= 1'b1;
24'h00a047: out <= 1'b1;
24'h00b047: out <= 1'b1;
24'h00c047: out <= 1'b1;
24'h00d047: out <= 1'b1;
24'h00e047: out <= 1'b1;
24'h00f047: out <= 1'b1;
24'h010047: out <= 1'b1;
24'h011047: out <= 1'b1;
24'h012047: out <= 1'b1;
24'h013047: out <= 1'b1;
24'h014047: out <= 1'b1;
24'h015047: out <= 1'b1;
24'h016047: out <= 1'b1;
24'h024047: out <= 1'b1;
24'h025047: out <= 1'b1;
24'h026047: out <= 1'b1;
24'h027047: out <= 1'b1;
24'h032047: out <= 1'b1;
24'h033047: out <= 1'b1;
24'h034047: out <= 1'b1;
24'h035047: out <= 1'b1;
24'h036047: out <= 1'b1;
24'h037047: out <= 1'b1;
24'h038047: out <= 1'b1;
24'h039047: out <= 1'b1;
24'h03a047: out <= 1'b1;
24'h03b047: out <= 1'b1;
24'h03c047: out <= 1'b1;
24'h03d047: out <= 1'b1;
24'h03e047: out <= 1'b1;
24'h03f047: out <= 1'b1;
24'h040047: out <= 1'b1;
24'h041047: out <= 1'b1;
24'h042047: out <= 1'b1;
24'h043047: out <= 1'b1;
24'h044047: out <= 1'b1;
24'h045047: out <= 1'b1;
24'h048047: out <= 1'b1;
24'h049047: out <= 1'b1;
24'h04a047: out <= 1'b1;
24'h04b047: out <= 1'b1;
24'h04c047: out <= 1'b1;
24'h04d047: out <= 1'b1;
24'h052047: out <= 1'b1;
24'h053047: out <= 1'b1;
24'h054047: out <= 1'b1;
24'h055047: out <= 1'b1;
24'h056047: out <= 1'b1;
24'h057047: out <= 1'b1;
24'h058047: out <= 1'b1;
24'h059047: out <= 1'b1;
24'h05a047: out <= 1'b1;
24'h05b047: out <= 1'b1;
default: out <= 1'b0;

endcase 
end
endmodule 