typedef logic [2:0] [63:0] vector;
typedef logic [63:0] fixed_real;
typedef logic [2:0] [7:0] color;

//javascript used to generate the long part
/*
function tobin(a){
	var str = Math.round(a * Math.pow(2,30));
	if(str < 0){
		var str1 = Math.abs(str).toString(2);
		var q = "1";
		for(var i = 0; i < 31-str1.length; i++){
			q += "0";
		}
		q += str1;
		return q;
	} else {
		return str.toString(2);
	}
}
var out = "always_ff @ (negedge Clk) begin\ncase (in)\n";
for(var i = 0; i <= 360; i++) {
		out += "9'd" + (i) + ": out <= 32'b"+tobin(Math.sin(i*Math.PI/180))+";    ";  //use cos for cos
		if(!(i % 3)){
			out += "\n";
		}
}
out += "endcase\nend\n";
console.log(out);
*/

module sin_lut(
	input logic Clk,
	input fixed_real angle,
	output fixed_real sin
);
fixed_real angle_fixed;
logic [8:0] in;
logic [15:0] out;
logic [14:0] out_fixed;


assign angle_fixed = angle[63]?angle+(64'd360 << 32):angle;

assign in = angle_fixed[40:32];
assign out_fixed = out[15]?(~out[14:0])+15'd1:out[14:0];
assign sin = {{31{out[15]}},out_fixed,18'd0};

always_ff @ (posedge Clk) begin
case (in)
9'd0: out <= 16'b0;    
9'd1: out <= 16'b100011110;    9'd2: out <= 16'b1000111100;    9'd3: out <= 16'b1101011001;    
9'd4: out <= 16'b10001110111;    9'd5: out <= 16'b10110010100;    9'd6: out <= 16'b11010110001;    
9'd7: out <= 16'b11111001101;    9'd8: out <= 16'b100011101000;    9'd9: out <= 16'b101000000011;    
9'd10: out <= 16'b101100011101;    9'd11: out <= 16'b110000110110;    9'd12: out <= 16'b110101001110;    
9'd13: out <= 16'b111001100110;    9'd14: out <= 16'b111101111100;    9'd15: out <= 16'b1000010010000;    
9'd16: out <= 16'b1000110100100;    9'd17: out <= 16'b1001010110110;    9'd18: out <= 16'b1001111000111;    
9'd19: out <= 16'b1010011010110;    9'd20: out <= 16'b1010111100100;    9'd21: out <= 16'b1011011110000;    
9'd22: out <= 16'b1011111111010;    9'd23: out <= 16'b1100100000010;    9'd24: out <= 16'b1101000001000;    
9'd25: out <= 16'b1101100001100;    9'd26: out <= 16'b1110000001110;    9'd27: out <= 16'b1110100001110;    
9'd28: out <= 16'b1111000001100;    9'd29: out <= 16'b1111100000111;    9'd30: out <= 16'b10000000000000;    
9'd31: out <= 16'b10000011110110;    9'd32: out <= 16'b10000111101010;    9'd33: out <= 16'b10001011011011;    
9'd34: out <= 16'b10001111001010;    9'd35: out <= 16'b10010010110101;    9'd36: out <= 16'b10010110011110;    
9'd37: out <= 16'b10011010000100;    9'd38: out <= 16'b10011101100111;    9'd39: out <= 16'b10100001000111;    
9'd40: out <= 16'b10100100100011;    9'd41: out <= 16'b10100111111101;    9'd42: out <= 16'b10101011010011;    
9'd43: out <= 16'b10101110100110;    9'd44: out <= 16'b10110001110101;    9'd45: out <= 16'b10110101000001;    
9'd46: out <= 16'b10111000001010;    9'd47: out <= 16'b10111011001110;    9'd48: out <= 16'b10111110010000;    
9'd49: out <= 16'b11000001001101;    9'd50: out <= 16'b11000100000111;    9'd51: out <= 16'b11000110111101;    
9'd52: out <= 16'b11001001101111;    9'd53: out <= 16'b11001100011101;    9'd54: out <= 16'b11001111000111;    
9'd55: out <= 16'b11010001101101;    9'd56: out <= 16'b11010100001111;    9'd57: out <= 16'b11010110101101;    
9'd58: out <= 16'b11011001000110;    9'd59: out <= 16'b11011011011100;    9'd60: out <= 16'b11011101101101;    
9'd61: out <= 16'b11011111111010;    9'd62: out <= 16'b11100010000010;    9'd63: out <= 16'b11100100000110;    
9'd64: out <= 16'b11100110000110;    9'd65: out <= 16'b11101000000001;    9'd66: out <= 16'b11101001111000;    
9'd67: out <= 16'b11101011101010;    9'd68: out <= 16'b11101101010111;    9'd69: out <= 16'b11101111000000;    
9'd70: out <= 16'b11110000100100;    9'd71: out <= 16'b11110010000011;    9'd72: out <= 16'b11110011011110;    
9'd73: out <= 16'b11110100110100;    9'd74: out <= 16'b11110110000101;    9'd75: out <= 16'b11110111010010;    
9'd76: out <= 16'b11111000011001;    9'd77: out <= 16'b11111001011100;    9'd78: out <= 16'b11111010011010;    
9'd79: out <= 16'b11111011010011;    9'd80: out <= 16'b11111100000111;    9'd81: out <= 16'b11111100110110;    
9'd82: out <= 16'b11111101100001;    9'd83: out <= 16'b11111110000110;    9'd84: out <= 16'b11111110100110;    
9'd85: out <= 16'b11111111000010;    9'd86: out <= 16'b11111111011000;    9'd87: out <= 16'b11111111101010;    
9'd88: out <= 16'b11111111110110;    9'd89: out <= 16'b11111111111110;    9'd90: out <= 16'b100000000000000;    
9'd91: out <= 16'b11111111111110;    9'd92: out <= 16'b11111111110110;    9'd93: out <= 16'b11111111101010;    
9'd94: out <= 16'b11111111011000;    9'd95: out <= 16'b11111111000010;    9'd96: out <= 16'b11111110100110;    
9'd97: out <= 16'b11111110000110;    9'd98: out <= 16'b11111101100001;    9'd99: out <= 16'b11111100110110;    
9'd100: out <= 16'b11111100000111;    9'd101: out <= 16'b11111011010011;    9'd102: out <= 16'b11111010011010;    
9'd103: out <= 16'b11111001011100;    9'd104: out <= 16'b11111000011001;    9'd105: out <= 16'b11110111010010;    
9'd106: out <= 16'b11110110000101;    9'd107: out <= 16'b11110100110100;    9'd108: out <= 16'b11110011011110;    
9'd109: out <= 16'b11110010000011;    9'd110: out <= 16'b11110000100100;    9'd111: out <= 16'b11101111000000;    
9'd112: out <= 16'b11101101010111;    9'd113: out <= 16'b11101011101010;    9'd114: out <= 16'b11101001111000;    
9'd115: out <= 16'b11101000000001;    9'd116: out <= 16'b11100110000110;    9'd117: out <= 16'b11100100000110;    
9'd118: out <= 16'b11100010000010;    9'd119: out <= 16'b11011111111010;    9'd120: out <= 16'b11011101101101;    
9'd121: out <= 16'b11011011011100;    9'd122: out <= 16'b11011001000110;    9'd123: out <= 16'b11010110101101;    
9'd124: out <= 16'b11010100001111;    9'd125: out <= 16'b11010001101101;    9'd126: out <= 16'b11001111000111;    
9'd127: out <= 16'b11001100011101;    9'd128: out <= 16'b11001001101111;    9'd129: out <= 16'b11000110111101;    
9'd130: out <= 16'b11000100000111;    9'd131: out <= 16'b11000001001101;    9'd132: out <= 16'b10111110010000;    
9'd133: out <= 16'b10111011001110;    9'd134: out <= 16'b10111000001010;    9'd135: out <= 16'b10110101000001;    
9'd136: out <= 16'b10110001110101;    9'd137: out <= 16'b10101110100110;    9'd138: out <= 16'b10101011010011;    
9'd139: out <= 16'b10100111111101;    9'd140: out <= 16'b10100100100011;    9'd141: out <= 16'b10100001000111;    
9'd142: out <= 16'b10011101100111;    9'd143: out <= 16'b10011010000100;    9'd144: out <= 16'b10010110011110;    
9'd145: out <= 16'b10010010110101;    9'd146: out <= 16'b10001111001010;    9'd147: out <= 16'b10001011011011;    
9'd148: out <= 16'b10000111101010;    9'd149: out <= 16'b10000011110110;    9'd150: out <= 16'b10000000000000;    
9'd151: out <= 16'b1111100000111;    9'd152: out <= 16'b1111000001100;    9'd153: out <= 16'b1110100001110;    
9'd154: out <= 16'b1110000001110;    9'd155: out <= 16'b1101100001100;    9'd156: out <= 16'b1101000001000;    
9'd157: out <= 16'b1100100000010;    9'd158: out <= 16'b1011111111010;    9'd159: out <= 16'b1011011110000;    
9'd160: out <= 16'b1010111100100;    9'd161: out <= 16'b1010011010110;    9'd162: out <= 16'b1001111000111;    
9'd163: out <= 16'b1001010110110;    9'd164: out <= 16'b1000110100100;    9'd165: out <= 16'b1000010010000;    
9'd166: out <= 16'b111101111100;    9'd167: out <= 16'b111001100110;    9'd168: out <= 16'b110101001110;    
9'd169: out <= 16'b110000110110;    9'd170: out <= 16'b101100011101;    9'd171: out <= 16'b101000000011;    
9'd172: out <= 16'b100011101000;    9'd173: out <= 16'b11111001101;    9'd174: out <= 16'b11010110001;    
9'd175: out <= 16'b10110010100;    9'd176: out <= 16'b10001110111;    9'd177: out <= 16'b1101011001;    
9'd178: out <= 16'b1000111100;    9'd179: out <= 16'b100011110;    9'd180: out <= 16'b0;    
9'd181: out <= 16'b1000000100011110;    9'd182: out <= 16'b1000001000111100;    9'd183: out <= 16'b1000001101011001;    
9'd184: out <= 16'b1000010001110111;    9'd185: out <= 16'b1000010110010100;    9'd186: out <= 16'b1000011010110001;    
9'd187: out <= 16'b1000011111001101;    9'd188: out <= 16'b1000100011101000;    9'd189: out <= 16'b1000101000000011;    
9'd190: out <= 16'b1000101100011101;    9'd191: out <= 16'b1000110000110110;    9'd192: out <= 16'b1000110101001110;    
9'd193: out <= 16'b1000111001100110;    9'd194: out <= 16'b1000111101111100;    9'd195: out <= 16'b1001000010010000;    
9'd196: out <= 16'b1001000110100100;    9'd197: out <= 16'b1001001010110110;    9'd198: out <= 16'b1001001111000111;    
9'd199: out <= 16'b1001010011010110;    9'd200: out <= 16'b1001010111100100;    9'd201: out <= 16'b1001011011110000;    
9'd202: out <= 16'b1001011111111010;    9'd203: out <= 16'b1001100100000010;    9'd204: out <= 16'b1001101000001000;    
9'd205: out <= 16'b1001101100001100;    9'd206: out <= 16'b1001110000001110;    9'd207: out <= 16'b1001110100001110;    
9'd208: out <= 16'b1001111000001100;    9'd209: out <= 16'b1001111100000111;    9'd210: out <= 16'b1010000000000000;    
9'd211: out <= 16'b1010000011110110;    9'd212: out <= 16'b1010000111101010;    9'd213: out <= 16'b1010001011011011;    
9'd214: out <= 16'b1010001111001010;    9'd215: out <= 16'b1010010010110101;    9'd216: out <= 16'b1010010110011110;    
9'd217: out <= 16'b1010011010000100;    9'd218: out <= 16'b1010011101100111;    9'd219: out <= 16'b1010100001000111;    
9'd220: out <= 16'b1010100100100011;    9'd221: out <= 16'b1010100111111101;    9'd222: out <= 16'b1010101011010011;    
9'd223: out <= 16'b1010101110100110;    9'd224: out <= 16'b1010110001110101;    9'd225: out <= 16'b1010110101000001;    
9'd226: out <= 16'b1010111000001010;    9'd227: out <= 16'b1010111011001110;    9'd228: out <= 16'b1010111110010000;    
9'd229: out <= 16'b1011000001001101;    9'd230: out <= 16'b1011000100000111;    9'd231: out <= 16'b1011000110111101;    
9'd232: out <= 16'b1011001001101111;    9'd233: out <= 16'b1011001100011101;    9'd234: out <= 16'b1011001111000111;    
9'd235: out <= 16'b1011010001101101;    9'd236: out <= 16'b1011010100001111;    9'd237: out <= 16'b1011010110101101;    
9'd238: out <= 16'b1011011001000110;    9'd239: out <= 16'b1011011011011100;    9'd240: out <= 16'b1011011101101101;    
9'd241: out <= 16'b1011011111111010;    9'd242: out <= 16'b1011100010000010;    9'd243: out <= 16'b1011100100000110;    
9'd244: out <= 16'b1011100110000110;    9'd245: out <= 16'b1011101000000001;    9'd246: out <= 16'b1011101001111000;    
9'd247: out <= 16'b1011101011101010;    9'd248: out <= 16'b1011101101010111;    9'd249: out <= 16'b1011101111000000;    
9'd250: out <= 16'b1011110000100100;    9'd251: out <= 16'b1011110010000011;    9'd252: out <= 16'b1011110011011110;    
9'd253: out <= 16'b1011110100110100;    9'd254: out <= 16'b1011110110000101;    9'd255: out <= 16'b1011110111010010;    
9'd256: out <= 16'b1011111000011001;    9'd257: out <= 16'b1011111001011100;    9'd258: out <= 16'b1011111010011010;    
9'd259: out <= 16'b1011111011010011;    9'd260: out <= 16'b1011111100000111;    9'd261: out <= 16'b1011111100110110;    
9'd262: out <= 16'b1011111101100001;    9'd263: out <= 16'b1011111110000110;    9'd264: out <= 16'b1011111110100110;    
9'd265: out <= 16'b1011111111000010;    9'd266: out <= 16'b1011111111011000;    9'd267: out <= 16'b1011111111101010;    
9'd268: out <= 16'b1011111111110110;    9'd269: out <= 16'b1011111111111110;    9'd270: out <= 16'b1100000000000000;    
9'd271: out <= 16'b1011111111111110;    9'd272: out <= 16'b1011111111110110;    9'd273: out <= 16'b1011111111101010;    
9'd274: out <= 16'b1011111111011000;    9'd275: out <= 16'b1011111111000010;    9'd276: out <= 16'b1011111110100110;    
9'd277: out <= 16'b1011111110000110;    9'd278: out <= 16'b1011111101100001;    9'd279: out <= 16'b1011111100110110;    
9'd280: out <= 16'b1011111100000111;    9'd281: out <= 16'b1011111011010011;    9'd282: out <= 16'b1011111010011010;    
9'd283: out <= 16'b1011111001011100;    9'd284: out <= 16'b1011111000011001;    9'd285: out <= 16'b1011110111010010;    
9'd286: out <= 16'b1011110110000101;    9'd287: out <= 16'b1011110100110100;    9'd288: out <= 16'b1011110011011110;    
9'd289: out <= 16'b1011110010000011;    9'd290: out <= 16'b1011110000100100;    9'd291: out <= 16'b1011101111000000;    
9'd292: out <= 16'b1011101101010111;    9'd293: out <= 16'b1011101011101010;    9'd294: out <= 16'b1011101001111000;    
9'd295: out <= 16'b1011101000000001;    9'd296: out <= 16'b1011100110000110;    9'd297: out <= 16'b1011100100000110;    
9'd298: out <= 16'b1011100010000010;    9'd299: out <= 16'b1011011111111010;    9'd300: out <= 16'b1011011101101101;    
9'd301: out <= 16'b1011011011011100;    9'd302: out <= 16'b1011011001000110;    9'd303: out <= 16'b1011010110101101;    
9'd304: out <= 16'b1011010100001111;    9'd305: out <= 16'b1011010001101101;    9'd306: out <= 16'b1011001111000111;    
9'd307: out <= 16'b1011001100011101;    9'd308: out <= 16'b1011001001101111;    9'd309: out <= 16'b1011000110111101;    
9'd310: out <= 16'b1011000100000111;    9'd311: out <= 16'b1011000001001101;    9'd312: out <= 16'b1010111110010000;    
9'd313: out <= 16'b1010111011001110;    9'd314: out <= 16'b1010111000001010;    9'd315: out <= 16'b1010110101000001;    
9'd316: out <= 16'b1010110001110101;    9'd317: out <= 16'b1010101110100110;    9'd318: out <= 16'b1010101011010011;    
9'd319: out <= 16'b1010100111111101;    9'd320: out <= 16'b1010100100100011;    9'd321: out <= 16'b1010100001000111;    
9'd322: out <= 16'b1010011101100111;    9'd323: out <= 16'b1010011010000100;    9'd324: out <= 16'b1010010110011110;    
9'd325: out <= 16'b1010010010110101;    9'd326: out <= 16'b1010001111001010;    9'd327: out <= 16'b1010001011011011;    
9'd328: out <= 16'b1010000111101010;    9'd329: out <= 16'b1010000011110110;    9'd330: out <= 16'b1010000000000000;    
9'd331: out <= 16'b1001111100000111;    9'd332: out <= 16'b1001111000001100;    9'd333: out <= 16'b1001110100001110;    
9'd334: out <= 16'b1001110000001110;    9'd335: out <= 16'b1001101100001100;    9'd336: out <= 16'b1001101000001000;    
9'd337: out <= 16'b1001100100000010;    9'd338: out <= 16'b1001011111111010;    9'd339: out <= 16'b1001011011110000;    
9'd340: out <= 16'b1001010111100100;    9'd341: out <= 16'b1001010011010110;    9'd342: out <= 16'b1001001111000111;    
9'd343: out <= 16'b1001001010110110;    9'd344: out <= 16'b1001000110100100;    9'd345: out <= 16'b1001000010010000;    
9'd346: out <= 16'b1000111101111100;    9'd347: out <= 16'b1000111001100110;    9'd348: out <= 16'b1000110101001110;    
9'd349: out <= 16'b1000110000110110;    9'd350: out <= 16'b1000101100011101;    9'd351: out <= 16'b1000101000000011;    
9'd352: out <= 16'b1000100011101000;    9'd353: out <= 16'b1000011111001101;    9'd354: out <= 16'b1000011010110001;    
9'd355: out <= 16'b1000010110010100;    9'd356: out <= 16'b1000010001110111;    9'd357: out <= 16'b1000001101011001;    
9'd358: out <= 16'b1000001000111100;    9'd359: out <= 16'b1000000100011110;    9'd360: out <= 16'b0;    
endcase
end


endmodule



module cos_lut(
	input logic Clk,
	input fixed_real angle,
	output fixed_real cos
);
fixed_real angle_fixed;
logic [8:0] in;
logic [15:0] out;
logic [14:0] out_fixed;


assign angle_fixed = angle[63]?angle+(64'd360 << 32):angle;

assign in = angle_fixed[40:32];
assign out_fixed = out[15]?(~out[14:0])+15'd1:out[14:0];
assign cos = {{31{out[15]}},out_fixed,18'd0};

always_ff @ (posedge Clk) begin
case (in)
9'd0: out <= 16'b100000000000000;    
9'd1: out <= 16'b11111111111110;    9'd2: out <= 16'b11111111110110;    9'd3: out <= 16'b11111111101010;    
9'd4: out <= 16'b11111111011000;    9'd5: out <= 16'b11111111000010;    9'd6: out <= 16'b11111110100110;    
9'd7: out <= 16'b11111110000110;    9'd8: out <= 16'b11111101100001;    9'd9: out <= 16'b11111100110110;    
9'd10: out <= 16'b11111100000111;    9'd11: out <= 16'b11111011010011;    9'd12: out <= 16'b11111010011010;    
9'd13: out <= 16'b11111001011100;    9'd14: out <= 16'b11111000011001;    9'd15: out <= 16'b11110111010010;    
9'd16: out <= 16'b11110110000101;    9'd17: out <= 16'b11110100110100;    9'd18: out <= 16'b11110011011110;    
9'd19: out <= 16'b11110010000011;    9'd20: out <= 16'b11110000100100;    9'd21: out <= 16'b11101111000000;    
9'd22: out <= 16'b11101101010111;    9'd23: out <= 16'b11101011101010;    9'd24: out <= 16'b11101001111000;    
9'd25: out <= 16'b11101000000001;    9'd26: out <= 16'b11100110000110;    9'd27: out <= 16'b11100100000110;    
9'd28: out <= 16'b11100010000010;    9'd29: out <= 16'b11011111111010;    9'd30: out <= 16'b11011101101101;    
9'd31: out <= 16'b11011011011100;    9'd32: out <= 16'b11011001000110;    9'd33: out <= 16'b11010110101101;    
9'd34: out <= 16'b11010100001111;    9'd35: out <= 16'b11010001101101;    9'd36: out <= 16'b11001111000111;    
9'd37: out <= 16'b11001100011101;    9'd38: out <= 16'b11001001101111;    9'd39: out <= 16'b11000110111101;    
9'd40: out <= 16'b11000100000111;    9'd41: out <= 16'b11000001001101;    9'd42: out <= 16'b10111110010000;    
9'd43: out <= 16'b10111011001110;    9'd44: out <= 16'b10111000001010;    9'd45: out <= 16'b10110101000001;    
9'd46: out <= 16'b10110001110101;    9'd47: out <= 16'b10101110100110;    9'd48: out <= 16'b10101011010011;    
9'd49: out <= 16'b10100111111101;    9'd50: out <= 16'b10100100100011;    9'd51: out <= 16'b10100001000111;    
9'd52: out <= 16'b10011101100111;    9'd53: out <= 16'b10011010000100;    9'd54: out <= 16'b10010110011110;    
9'd55: out <= 16'b10010010110101;    9'd56: out <= 16'b10001111001010;    9'd57: out <= 16'b10001011011011;    
9'd58: out <= 16'b10000111101010;    9'd59: out <= 16'b10000011110110;    9'd60: out <= 16'b10000000000000;    
9'd61: out <= 16'b1111100000111;    9'd62: out <= 16'b1111000001100;    9'd63: out <= 16'b1110100001110;    
9'd64: out <= 16'b1110000001110;    9'd65: out <= 16'b1101100001100;    9'd66: out <= 16'b1101000001000;    
9'd67: out <= 16'b1100100000010;    9'd68: out <= 16'b1011111111010;    9'd69: out <= 16'b1011011110000;    
9'd70: out <= 16'b1010111100100;    9'd71: out <= 16'b1010011010110;    9'd72: out <= 16'b1001111000111;    
9'd73: out <= 16'b1001010110110;    9'd74: out <= 16'b1000110100100;    9'd75: out <= 16'b1000010010000;    
9'd76: out <= 16'b111101111100;    9'd77: out <= 16'b111001100110;    9'd78: out <= 16'b110101001110;    
9'd79: out <= 16'b110000110110;    9'd80: out <= 16'b101100011101;    9'd81: out <= 16'b101000000011;    
9'd82: out <= 16'b100011101000;    9'd83: out <= 16'b11111001101;    9'd84: out <= 16'b11010110001;    
9'd85: out <= 16'b10110010100;    9'd86: out <= 16'b10001110111;    9'd87: out <= 16'b1101011001;    
9'd88: out <= 16'b1000111100;    9'd89: out <= 16'b100011110;    9'd90: out <= 16'b0;    
9'd91: out <= 16'b1000000100011110;    9'd92: out <= 16'b1000001000111100;    9'd93: out <= 16'b1000001101011001;    
9'd94: out <= 16'b1000010001110111;    9'd95: out <= 16'b1000010110010100;    9'd96: out <= 16'b1000011010110001;    
9'd97: out <= 16'b1000011111001101;    9'd98: out <= 16'b1000100011101000;    9'd99: out <= 16'b1000101000000011;    
9'd100: out <= 16'b1000101100011101;    9'd101: out <= 16'b1000110000110110;    9'd102: out <= 16'b1000110101001110;    
9'd103: out <= 16'b1000111001100110;    9'd104: out <= 16'b1000111101111100;    9'd105: out <= 16'b1001000010010000;    
9'd106: out <= 16'b1001000110100100;    9'd107: out <= 16'b1001001010110110;    9'd108: out <= 16'b1001001111000111;    
9'd109: out <= 16'b1001010011010110;    9'd110: out <= 16'b1001010111100100;    9'd111: out <= 16'b1001011011110000;    
9'd112: out <= 16'b1001011111111010;    9'd113: out <= 16'b1001100100000010;    9'd114: out <= 16'b1001101000001000;    
9'd115: out <= 16'b1001101100001100;    9'd116: out <= 16'b1001110000001110;    9'd117: out <= 16'b1001110100001110;    
9'd118: out <= 16'b1001111000001100;    9'd119: out <= 16'b1001111100000111;    9'd120: out <= 16'b1010000000000000;    
9'd121: out <= 16'b1010000011110110;    9'd122: out <= 16'b1010000111101010;    9'd123: out <= 16'b1010001011011011;    
9'd124: out <= 16'b1010001111001010;    9'd125: out <= 16'b1010010010110101;    9'd126: out <= 16'b1010010110011110;    
9'd127: out <= 16'b1010011010000100;    9'd128: out <= 16'b1010011101100111;    9'd129: out <= 16'b1010100001000111;    
9'd130: out <= 16'b1010100100100011;    9'd131: out <= 16'b1010100111111101;    9'd132: out <= 16'b1010101011010011;    
9'd133: out <= 16'b1010101110100110;    9'd134: out <= 16'b1010110001110101;    9'd135: out <= 16'b1010110101000001;    
9'd136: out <= 16'b1010111000001010;    9'd137: out <= 16'b1010111011001110;    9'd138: out <= 16'b1010111110010000;    
9'd139: out <= 16'b1011000001001101;    9'd140: out <= 16'b1011000100000111;    9'd141: out <= 16'b1011000110111101;    
9'd142: out <= 16'b1011001001101111;    9'd143: out <= 16'b1011001100011101;    9'd144: out <= 16'b1011001111000111;    
9'd145: out <= 16'b1011010001101101;    9'd146: out <= 16'b1011010100001111;    9'd147: out <= 16'b1011010110101101;    
9'd148: out <= 16'b1011011001000110;    9'd149: out <= 16'b1011011011011100;    9'd150: out <= 16'b1011011101101101;    
9'd151: out <= 16'b1011011111111010;    9'd152: out <= 16'b1011100010000010;    9'd153: out <= 16'b1011100100000110;    
9'd154: out <= 16'b1011100110000110;    9'd155: out <= 16'b1011101000000001;    9'd156: out <= 16'b1011101001111000;    
9'd157: out <= 16'b1011101011101010;    9'd158: out <= 16'b1011101101010111;    9'd159: out <= 16'b1011101111000000;    
9'd160: out <= 16'b1011110000100100;    9'd161: out <= 16'b1011110010000011;    9'd162: out <= 16'b1011110011011110;    
9'd163: out <= 16'b1011110100110100;    9'd164: out <= 16'b1011110110000101;    9'd165: out <= 16'b1011110111010010;    
9'd166: out <= 16'b1011111000011001;    9'd167: out <= 16'b1011111001011100;    9'd168: out <= 16'b1011111010011010;    
9'd169: out <= 16'b1011111011010011;    9'd170: out <= 16'b1011111100000111;    9'd171: out <= 16'b1011111100110110;    
9'd172: out <= 16'b1011111101100001;    9'd173: out <= 16'b1011111110000110;    9'd174: out <= 16'b1011111110100110;    
9'd175: out <= 16'b1011111111000010;    9'd176: out <= 16'b1011111111011000;    9'd177: out <= 16'b1011111111101010;    
9'd178: out <= 16'b1011111111110110;    9'd179: out <= 16'b1011111111111110;    9'd180: out <= 16'b1100000000000000;    
9'd181: out <= 16'b1011111111111110;    9'd182: out <= 16'b1011111111110110;    9'd183: out <= 16'b1011111111101010;    
9'd184: out <= 16'b1011111111011000;    9'd185: out <= 16'b1011111111000010;    9'd186: out <= 16'b1011111110100110;    
9'd187: out <= 16'b1011111110000110;    9'd188: out <= 16'b1011111101100001;    9'd189: out <= 16'b1011111100110110;    
9'd190: out <= 16'b1011111100000111;    9'd191: out <= 16'b1011111011010011;    9'd192: out <= 16'b1011111010011010;    
9'd193: out <= 16'b1011111001011100;    9'd194: out <= 16'b1011111000011001;    9'd195: out <= 16'b1011110111010010;    
9'd196: out <= 16'b1011110110000101;    9'd197: out <= 16'b1011110100110100;    9'd198: out <= 16'b1011110011011110;    
9'd199: out <= 16'b1011110010000011;    9'd200: out <= 16'b1011110000100100;    9'd201: out <= 16'b1011101111000000;    
9'd202: out <= 16'b1011101101010111;    9'd203: out <= 16'b1011101011101010;    9'd204: out <= 16'b1011101001111000;    
9'd205: out <= 16'b1011101000000001;    9'd206: out <= 16'b1011100110000110;    9'd207: out <= 16'b1011100100000110;    
9'd208: out <= 16'b1011100010000010;    9'd209: out <= 16'b1011011111111010;    9'd210: out <= 16'b1011011101101101;    
9'd211: out <= 16'b1011011011011100;    9'd212: out <= 16'b1011011001000110;    9'd213: out <= 16'b1011010110101101;    
9'd214: out <= 16'b1011010100001111;    9'd215: out <= 16'b1011010001101101;    9'd216: out <= 16'b1011001111000111;    
9'd217: out <= 16'b1011001100011101;    9'd218: out <= 16'b1011001001101111;    9'd219: out <= 16'b1011000110111101;    
9'd220: out <= 16'b1011000100000111;    9'd221: out <= 16'b1011000001001101;    9'd222: out <= 16'b1010111110010000;    
9'd223: out <= 16'b1010111011001110;    9'd224: out <= 16'b1010111000001010;    9'd225: out <= 16'b1010110101000001;    
9'd226: out <= 16'b1010110001110101;    9'd227: out <= 16'b1010101110100110;    9'd228: out <= 16'b1010101011010011;    
9'd229: out <= 16'b1010100111111101;    9'd230: out <= 16'b1010100100100011;    9'd231: out <= 16'b1010100001000111;    
9'd232: out <= 16'b1010011101100111;    9'd233: out <= 16'b1010011010000100;    9'd234: out <= 16'b1010010110011110;    
9'd235: out <= 16'b1010010010110101;    9'd236: out <= 16'b1010001111001010;    9'd237: out <= 16'b1010001011011011;    
9'd238: out <= 16'b1010000111101010;    9'd239: out <= 16'b1010000011110110;    9'd240: out <= 16'b1010000000000000;    
9'd241: out <= 16'b1001111100000111;    9'd242: out <= 16'b1001111000001100;    9'd243: out <= 16'b1001110100001110;    
9'd244: out <= 16'b1001110000001110;    9'd245: out <= 16'b1001101100001100;    9'd246: out <= 16'b1001101000001000;    
9'd247: out <= 16'b1001100100000010;    9'd248: out <= 16'b1001011111111010;    9'd249: out <= 16'b1001011011110000;    
9'd250: out <= 16'b1001010111100100;    9'd251: out <= 16'b1001010011010110;    9'd252: out <= 16'b1001001111000111;    
9'd253: out <= 16'b1001001010110110;    9'd254: out <= 16'b1001000110100100;    9'd255: out <= 16'b1001000010010000;    
9'd256: out <= 16'b1000111101111100;    9'd257: out <= 16'b1000111001100110;    9'd258: out <= 16'b1000110101001110;    
9'd259: out <= 16'b1000110000110110;    9'd260: out <= 16'b1000101100011101;    9'd261: out <= 16'b1000101000000011;    
9'd262: out <= 16'b1000100011101000;    9'd263: out <= 16'b1000011111001101;    9'd264: out <= 16'b1000011010110001;    
9'd265: out <= 16'b1000010110010100;    9'd266: out <= 16'b1000010001110111;    9'd267: out <= 16'b1000001101011001;    
9'd268: out <= 16'b1000001000111100;    9'd269: out <= 16'b1000000100011110;    9'd270: out <= 16'b0;    
9'd271: out <= 16'b100011110;    9'd272: out <= 16'b1000111100;    9'd273: out <= 16'b1101011001;    
9'd274: out <= 16'b10001110111;    9'd275: out <= 16'b10110010100;    9'd276: out <= 16'b11010110001;    
9'd277: out <= 16'b11111001101;    9'd278: out <= 16'b100011101000;    9'd279: out <= 16'b101000000011;    
9'd280: out <= 16'b101100011101;    9'd281: out <= 16'b110000110110;    9'd282: out <= 16'b110101001110;    
9'd283: out <= 16'b111001100110;    9'd284: out <= 16'b111101111100;    9'd285: out <= 16'b1000010010000;    
9'd286: out <= 16'b1000110100100;    9'd287: out <= 16'b1001010110110;    9'd288: out <= 16'b1001111000111;    
9'd289: out <= 16'b1010011010110;    9'd290: out <= 16'b1010111100100;    9'd291: out <= 16'b1011011110000;    
9'd292: out <= 16'b1011111111010;    9'd293: out <= 16'b1100100000010;    9'd294: out <= 16'b1101000001000;    
9'd295: out <= 16'b1101100001100;    9'd296: out <= 16'b1110000001110;    9'd297: out <= 16'b1110100001110;    
9'd298: out <= 16'b1111000001100;    9'd299: out <= 16'b1111100000111;    9'd300: out <= 16'b10000000000000;    
9'd301: out <= 16'b10000011110110;    9'd302: out <= 16'b10000111101010;    9'd303: out <= 16'b10001011011011;    
9'd304: out <= 16'b10001111001010;    9'd305: out <= 16'b10010010110101;    9'd306: out <= 16'b10010110011110;    
9'd307: out <= 16'b10011010000100;    9'd308: out <= 16'b10011101100111;    9'd309: out <= 16'b10100001000111;    
9'd310: out <= 16'b10100100100011;    9'd311: out <= 16'b10100111111101;    9'd312: out <= 16'b10101011010011;    
9'd313: out <= 16'b10101110100110;    9'd314: out <= 16'b10110001110101;    9'd315: out <= 16'b10110101000001;    
9'd316: out <= 16'b10111000001010;    9'd317: out <= 16'b10111011001110;    9'd318: out <= 16'b10111110010000;    
9'd319: out <= 16'b11000001001101;    9'd320: out <= 16'b11000100000111;    9'd321: out <= 16'b11000110111101;    
9'd322: out <= 16'b11001001101111;    9'd323: out <= 16'b11001100011101;    9'd324: out <= 16'b11001111000111;    
9'd325: out <= 16'b11010001101101;    9'd326: out <= 16'b11010100001111;    9'd327: out <= 16'b11010110101101;    
9'd328: out <= 16'b11011001000110;    9'd329: out <= 16'b11011011011100;    9'd330: out <= 16'b11011101101101;    
9'd331: out <= 16'b11011111111010;    9'd332: out <= 16'b11100010000010;    9'd333: out <= 16'b11100100000110;    
9'd334: out <= 16'b11100110000110;    9'd335: out <= 16'b11101000000001;    9'd336: out <= 16'b11101001111000;    
9'd337: out <= 16'b11101011101010;    9'd338: out <= 16'b11101101010111;    9'd339: out <= 16'b11101111000000;    
9'd340: out <= 16'b11110000100100;    9'd341: out <= 16'b11110010000011;    9'd342: out <= 16'b11110011011110;    
9'd343: out <= 16'b11110100110100;    9'd344: out <= 16'b11110110000101;    9'd345: out <= 16'b11110111010010;    
9'd346: out <= 16'b11111000011001;    9'd347: out <= 16'b11111001011100;    9'd348: out <= 16'b11111010011010;    
9'd349: out <= 16'b11111011010011;    9'd350: out <= 16'b11111100000111;    9'd351: out <= 16'b11111100110110;    
9'd352: out <= 16'b11111101100001;    9'd353: out <= 16'b11111110000110;    9'd354: out <= 16'b11111110100110;    
9'd355: out <= 16'b11111111000010;    9'd356: out <= 16'b11111111011000;    9'd357: out <= 16'b11111111101010;    
9'd358: out <= 16'b11111111110110;    9'd359: out <= 16'b11111111111110;    9'd360: out <= 16'b100000000000000;    
endcase
end

endmodule

module ray_lut(
	input logic Clk,
	input fixed_real theta, phi,
	output vector ray
);

fixed_real cosTheta, sinTheta, sinPhi, cosPhi,x,y,z;

sin_lut s0(.*,.angle(theta),.sin(sinTheta));
sin_lut s1(.*,.angle(phi),.sin(sinPhi));
cos_lut c0(.*,.angle(theta),.cos(cosTheta));
cos_lut c1(.*,.angle(phi),.cos(cosPhi));

mult_real m0(.a(sinTheta),.b(sinPhi),.c(y));
mult_real m1(.a(sinTheta),.b(cosPhi),.c(z));

assign x = cosTheta;

assign ray = {z,y,x};

endmodule
