module pauselut (input [23:0] in, input Clk, output out);


always_ff @ (posedge Clk) begin
case (in)


24'h005029: out <= 1'b1;
24'h006029: out <= 1'b1;
24'h007029: out <= 1'b1;
24'h008029: out <= 1'b1;
24'h009029: out <= 1'b1;
24'h00a029: out <= 1'b1;
24'h00b029: out <= 1'b1;
24'h017029: out <= 1'b1;
24'h018029: out <= 1'b1;
24'h019029: out <= 1'b1;
24'h020029: out <= 1'b1;
24'h021029: out <= 1'b1;
24'h02a029: out <= 1'b1;
24'h02b029: out <= 1'b1;
24'h034029: out <= 1'b1;
24'h035029: out <= 1'b1;
24'h036029: out <= 1'b1;
24'h037029: out <= 1'b1;
24'h038029: out <= 1'b1;
24'h039029: out <= 1'b1;
24'h03a029: out <= 1'b1;
24'h03e029: out <= 1'b1;
24'h03f029: out <= 1'b1;
24'h040029: out <= 1'b1;
24'h041029: out <= 1'b1;
24'h042029: out <= 1'b1;
24'h043029: out <= 1'b1;
24'h044029: out <= 1'b1;
24'h045029: out <= 1'b1;
24'h046029: out <= 1'b1;
24'h047029: out <= 1'b1;
24'h048029: out <= 1'b1;
24'h04c029: out <= 1'b1;
24'h04d029: out <= 1'b1;
24'h04e029: out <= 1'b1;
24'h04f029: out <= 1'b1;
24'h00502a: out <= 1'b1;
24'h00602a: out <= 1'b1;
24'h00702a: out <= 1'b1;
24'h00802a: out <= 1'b1;
24'h00902a: out <= 1'b1;
24'h00a02a: out <= 1'b1;
24'h00b02a: out <= 1'b1;
24'h00c02a: out <= 1'b1;
24'h01702a: out <= 1'b1;
24'h01802a: out <= 1'b1;
24'h01902a: out <= 1'b1;
24'h02002a: out <= 1'b1;
24'h02102a: out <= 1'b1;
24'h02a02a: out <= 1'b1;
24'h02b02a: out <= 1'b1;
24'h03302a: out <= 1'b1;
24'h03402a: out <= 1'b1;
24'h03502a: out <= 1'b1;
24'h03602a: out <= 1'b1;
24'h03702a: out <= 1'b1;
24'h03802a: out <= 1'b1;
24'h03902a: out <= 1'b1;
24'h03a02a: out <= 1'b1;
24'h03e02a: out <= 1'b1;
24'h03f02a: out <= 1'b1;
24'h04002a: out <= 1'b1;
24'h04102a: out <= 1'b1;
24'h04202a: out <= 1'b1;
24'h04302a: out <= 1'b1;
24'h04402a: out <= 1'b1;
24'h04502a: out <= 1'b1;
24'h04602a: out <= 1'b1;
24'h04702a: out <= 1'b1;
24'h04802a: out <= 1'b1;
24'h04c02a: out <= 1'b1;
24'h04d02a: out <= 1'b1;
24'h04e02a: out <= 1'b1;
24'h04f02a: out <= 1'b1;
24'h05002a: out <= 1'b1;
24'h05102a: out <= 1'b1;
24'h00502b: out <= 1'b1;
24'h00602b: out <= 1'b1;
24'h00902b: out <= 1'b1;
24'h00a02b: out <= 1'b1;
24'h00b02b: out <= 1'b1;
24'h00c02b: out <= 1'b1;
24'h00d02b: out <= 1'b1;
24'h01602b: out <= 1'b1;
24'h01702b: out <= 1'b1;
24'h01802b: out <= 1'b1;
24'h01902b: out <= 1'b1;
24'h01a02b: out <= 1'b1;
24'h02002b: out <= 1'b1;
24'h02102b: out <= 1'b1;
24'h02a02b: out <= 1'b1;
24'h02b02b: out <= 1'b1;
24'h03202b: out <= 1'b1;
24'h03302b: out <= 1'b1;
24'h03402b: out <= 1'b1;
24'h03502b: out <= 1'b1;
24'h03602b: out <= 1'b1;
24'h03e02b: out <= 1'b1;
24'h03f02b: out <= 1'b1;
24'h04c02b: out <= 1'b1;
24'h04d02b: out <= 1'b1;
24'h04e02b: out <= 1'b1;
24'h04f02b: out <= 1'b1;
24'h05002b: out <= 1'b1;
24'h05102b: out <= 1'b1;
24'h05202b: out <= 1'b1;
24'h05302b: out <= 1'b1;
24'h00502c: out <= 1'b1;
24'h00602c: out <= 1'b1;
24'h00b02c: out <= 1'b1;
24'h00c02c: out <= 1'b1;
24'h00d02c: out <= 1'b1;
24'h01502c: out <= 1'b1;
24'h01602c: out <= 1'b1;
24'h01702c: out <= 1'b1;
24'h01802c: out <= 1'b1;
24'h01902c: out <= 1'b1;
24'h01a02c: out <= 1'b1;
24'h02002c: out <= 1'b1;
24'h02102c: out <= 1'b1;
24'h02a02c: out <= 1'b1;
24'h02b02c: out <= 1'b1;
24'h03102c: out <= 1'b1;
24'h03202c: out <= 1'b1;
24'h03302c: out <= 1'b1;
24'h03e02c: out <= 1'b1;
24'h03f02c: out <= 1'b1;
24'h04c02c: out <= 1'b1;
24'h04d02c: out <= 1'b1;
24'h05002c: out <= 1'b1;
24'h05102c: out <= 1'b1;
24'h05202c: out <= 1'b1;
24'h05302c: out <= 1'b1;
24'h05402c: out <= 1'b1;
24'h00502d: out <= 1'b1;
24'h00602d: out <= 1'b1;
24'h00c02d: out <= 1'b1;
24'h00d02d: out <= 1'b1;
24'h01502d: out <= 1'b1;
24'h01602d: out <= 1'b1;
24'h01702d: out <= 1'b1;
24'h01802d: out <= 1'b1;
24'h01902d: out <= 1'b1;
24'h01a02d: out <= 1'b1;
24'h02002d: out <= 1'b1;
24'h02102d: out <= 1'b1;
24'h02a02d: out <= 1'b1;
24'h02b02d: out <= 1'b1;
24'h03102d: out <= 1'b1;
24'h03202d: out <= 1'b1;
24'h03302d: out <= 1'b1;
24'h03e02d: out <= 1'b1;
24'h03f02d: out <= 1'b1;
24'h04c02d: out <= 1'b1;
24'h04d02d: out <= 1'b1;
24'h05202d: out <= 1'b1;
24'h05302d: out <= 1'b1;
24'h05402d: out <= 1'b1;
24'h05502d: out <= 1'b1;
24'h00502e: out <= 1'b1;
24'h00602e: out <= 1'b1;
24'h00b02e: out <= 1'b1;
24'h00c02e: out <= 1'b1;
24'h00d02e: out <= 1'b1;
24'h01402e: out <= 1'b1;
24'h01502e: out <= 1'b1;
24'h01602e: out <= 1'b1;
24'h01702e: out <= 1'b1;
24'h01802e: out <= 1'b1;
24'h01902e: out <= 1'b1;
24'h01a02e: out <= 1'b1;
24'h02002e: out <= 1'b1;
24'h02102e: out <= 1'b1;
24'h02a02e: out <= 1'b1;
24'h02b02e: out <= 1'b1;
24'h03102e: out <= 1'b1;
24'h03202e: out <= 1'b1;
24'h03302e: out <= 1'b1;
24'h03e02e: out <= 1'b1;
24'h03f02e: out <= 1'b1;
24'h04c02e: out <= 1'b1;
24'h04d02e: out <= 1'b1;
24'h05402e: out <= 1'b1;
24'h05502e: out <= 1'b1;
24'h05602e: out <= 1'b1;
24'h00502f: out <= 1'b1;
24'h00602f: out <= 1'b1;
24'h00b02f: out <= 1'b1;
24'h00c02f: out <= 1'b1;
24'h00d02f: out <= 1'b1;
24'h01302f: out <= 1'b1;
24'h01402f: out <= 1'b1;
24'h01502f: out <= 1'b1;
24'h01602f: out <= 1'b1;
24'h01702f: out <= 1'b1;
24'h01902f: out <= 1'b1;
24'h01a02f: out <= 1'b1;
24'h02002f: out <= 1'b1;
24'h02102f: out <= 1'b1;
24'h02902f: out <= 1'b1;
24'h02a02f: out <= 1'b1;
24'h02b02f: out <= 1'b1;
24'h03102f: out <= 1'b1;
24'h03202f: out <= 1'b1;
24'h03302f: out <= 1'b1;
24'h03402f: out <= 1'b1;
24'h03502f: out <= 1'b1;
24'h03e02f: out <= 1'b1;
24'h03f02f: out <= 1'b1;
24'h04002f: out <= 1'b1;
24'h04102f: out <= 1'b1;
24'h04202f: out <= 1'b1;
24'h04302f: out <= 1'b1;
24'h04402f: out <= 1'b1;
24'h04502f: out <= 1'b1;
24'h04602f: out <= 1'b1;
24'h04702f: out <= 1'b1;
24'h04c02f: out <= 1'b1;
24'h04d02f: out <= 1'b1;
24'h05502f: out <= 1'b1;
24'h05602f: out <= 1'b1;
24'h05702f: out <= 1'b1;
24'h005030: out <= 1'b1;
24'h006030: out <= 1'b1;
24'h007030: out <= 1'b1;
24'h009030: out <= 1'b1;
24'h00a030: out <= 1'b1;
24'h00b030: out <= 1'b1;
24'h00c030: out <= 1'b1;
24'h00d030: out <= 1'b1;
24'h013030: out <= 1'b1;
24'h014030: out <= 1'b1;
24'h015030: out <= 1'b1;
24'h016030: out <= 1'b1;
24'h019030: out <= 1'b1;
24'h01a030: out <= 1'b1;
24'h01b030: out <= 1'b1;
24'h020030: out <= 1'b1;
24'h021030: out <= 1'b1;
24'h029030: out <= 1'b1;
24'h02a030: out <= 1'b1;
24'h02b030: out <= 1'b1;
24'h031030: out <= 1'b1;
24'h032030: out <= 1'b1;
24'h033030: out <= 1'b1;
24'h034030: out <= 1'b1;
24'h035030: out <= 1'b1;
24'h036030: out <= 1'b1;
24'h037030: out <= 1'b1;
24'h038030: out <= 1'b1;
24'h039030: out <= 1'b1;
24'h03e030: out <= 1'b1;
24'h03f030: out <= 1'b1;
24'h040030: out <= 1'b1;
24'h041030: out <= 1'b1;
24'h042030: out <= 1'b1;
24'h043030: out <= 1'b1;
24'h044030: out <= 1'b1;
24'h045030: out <= 1'b1;
24'h046030: out <= 1'b1;
24'h047030: out <= 1'b1;
24'h04c030: out <= 1'b1;
24'h04d030: out <= 1'b1;
24'h055030: out <= 1'b1;
24'h056030: out <= 1'b1;
24'h057030: out <= 1'b1;
24'h005031: out <= 1'b1;
24'h006031: out <= 1'b1;
24'h007031: out <= 1'b1;
24'h008031: out <= 1'b1;
24'h009031: out <= 1'b1;
24'h00a031: out <= 1'b1;
24'h00b031: out <= 1'b1;
24'h00c031: out <= 1'b1;
24'h012031: out <= 1'b1;
24'h013031: out <= 1'b1;
24'h014031: out <= 1'b1;
24'h015031: out <= 1'b1;
24'h016031: out <= 1'b1;
24'h017031: out <= 1'b1;
24'h018031: out <= 1'b1;
24'h019031: out <= 1'b1;
24'h01a031: out <= 1'b1;
24'h01b031: out <= 1'b1;
24'h020031: out <= 1'b1;
24'h021031: out <= 1'b1;
24'h029031: out <= 1'b1;
24'h02a031: out <= 1'b1;
24'h02b031: out <= 1'b1;
24'h032031: out <= 1'b1;
24'h033031: out <= 1'b1;
24'h034031: out <= 1'b1;
24'h035031: out <= 1'b1;
24'h036031: out <= 1'b1;
24'h037031: out <= 1'b1;
24'h038031: out <= 1'b1;
24'h039031: out <= 1'b1;
24'h03a031: out <= 1'b1;
24'h03e031: out <= 1'b1;
24'h03f031: out <= 1'b1;
24'h040031: out <= 1'b1;
24'h041031: out <= 1'b1;
24'h042031: out <= 1'b1;
24'h043031: out <= 1'b1;
24'h044031: out <= 1'b1;
24'h045031: out <= 1'b1;
24'h046031: out <= 1'b1;
24'h04c031: out <= 1'b1;
24'h04d031: out <= 1'b1;
24'h055031: out <= 1'b1;
24'h056031: out <= 1'b1;
24'h057031: out <= 1'b1;
24'h005032: out <= 1'b1;
24'h006032: out <= 1'b1;
24'h007032: out <= 1'b1;
24'h008032: out <= 1'b1;
24'h009032: out <= 1'b1;
24'h00a032: out <= 1'b1;
24'h00b032: out <= 1'b1;
24'h011032: out <= 1'b1;
24'h012032: out <= 1'b1;
24'h013032: out <= 1'b1;
24'h014032: out <= 1'b1;
24'h015032: out <= 1'b1;
24'h016032: out <= 1'b1;
24'h017032: out <= 1'b1;
24'h018032: out <= 1'b1;
24'h019032: out <= 1'b1;
24'h01a032: out <= 1'b1;
24'h01b032: out <= 1'b1;
24'h020032: out <= 1'b1;
24'h021032: out <= 1'b1;
24'h022032: out <= 1'b1;
24'h029032: out <= 1'b1;
24'h02a032: out <= 1'b1;
24'h02b032: out <= 1'b1;
24'h036032: out <= 1'b1;
24'h037032: out <= 1'b1;
24'h038032: out <= 1'b1;
24'h039032: out <= 1'b1;
24'h03a032: out <= 1'b1;
24'h03b032: out <= 1'b1;
24'h03e032: out <= 1'b1;
24'h03f032: out <= 1'b1;
24'h04c032: out <= 1'b1;
24'h04d032: out <= 1'b1;
24'h056032: out <= 1'b1;
24'h057032: out <= 1'b1;
24'h005033: out <= 1'b1;
24'h006033: out <= 1'b1;
24'h011033: out <= 1'b1;
24'h012033: out <= 1'b1;
24'h013033: out <= 1'b1;
24'h014033: out <= 1'b1;
24'h015033: out <= 1'b1;
24'h016033: out <= 1'b1;
24'h017033: out <= 1'b1;
24'h018033: out <= 1'b1;
24'h019033: out <= 1'b1;
24'h01a033: out <= 1'b1;
24'h01b033: out <= 1'b1;
24'h020033: out <= 1'b1;
24'h021033: out <= 1'b1;
24'h022033: out <= 1'b1;
24'h029033: out <= 1'b1;
24'h02a033: out <= 1'b1;
24'h02b033: out <= 1'b1;
24'h039033: out <= 1'b1;
24'h03a033: out <= 1'b1;
24'h03b033: out <= 1'b1;
24'h03e033: out <= 1'b1;
24'h03f033: out <= 1'b1;
24'h04c033: out <= 1'b1;
24'h04d033: out <= 1'b1;
24'h055033: out <= 1'b1;
24'h056033: out <= 1'b1;
24'h057033: out <= 1'b1;
24'h005034: out <= 1'b1;
24'h006034: out <= 1'b1;
24'h011034: out <= 1'b1;
24'h012034: out <= 1'b1;
24'h013034: out <= 1'b1;
24'h014034: out <= 1'b1;
24'h01a034: out <= 1'b1;
24'h01b034: out <= 1'b1;
24'h020034: out <= 1'b1;
24'h021034: out <= 1'b1;
24'h022034: out <= 1'b1;
24'h028034: out <= 1'b1;
24'h029034: out <= 1'b1;
24'h02a034: out <= 1'b1;
24'h02b034: out <= 1'b1;
24'h03a034: out <= 1'b1;
24'h03b034: out <= 1'b1;
24'h03e034: out <= 1'b1;
24'h03f034: out <= 1'b1;
24'h04c034: out <= 1'b1;
24'h04d034: out <= 1'b1;
24'h055034: out <= 1'b1;
24'h056034: out <= 1'b1;
24'h057034: out <= 1'b1;
24'h005035: out <= 1'b1;
24'h006035: out <= 1'b1;
24'h010035: out <= 1'b1;
24'h011035: out <= 1'b1;
24'h012035: out <= 1'b1;
24'h013035: out <= 1'b1;
24'h01a035: out <= 1'b1;
24'h01b035: out <= 1'b1;
24'h01c035: out <= 1'b1;
24'h020035: out <= 1'b1;
24'h021035: out <= 1'b1;
24'h022035: out <= 1'b1;
24'h023035: out <= 1'b1;
24'h028035: out <= 1'b1;
24'h029035: out <= 1'b1;
24'h02a035: out <= 1'b1;
24'h039035: out <= 1'b1;
24'h03a035: out <= 1'b1;
24'h03b035: out <= 1'b1;
24'h03e035: out <= 1'b1;
24'h03f035: out <= 1'b1;
24'h04c035: out <= 1'b1;
24'h04d035: out <= 1'b1;
24'h054035: out <= 1'b1;
24'h055035: out <= 1'b1;
24'h056035: out <= 1'b1;
24'h057035: out <= 1'b1;
24'h005036: out <= 1'b1;
24'h006036: out <= 1'b1;
24'h010036: out <= 1'b1;
24'h011036: out <= 1'b1;
24'h012036: out <= 1'b1;
24'h013036: out <= 1'b1;
24'h01a036: out <= 1'b1;
24'h01b036: out <= 1'b1;
24'h01c036: out <= 1'b1;
24'h021036: out <= 1'b1;
24'h022036: out <= 1'b1;
24'h023036: out <= 1'b1;
24'h024036: out <= 1'b1;
24'h025036: out <= 1'b1;
24'h026036: out <= 1'b1;
24'h027036: out <= 1'b1;
24'h028036: out <= 1'b1;
24'h029036: out <= 1'b1;
24'h02a036: out <= 1'b1;
24'h030036: out <= 1'b1;
24'h031036: out <= 1'b1;
24'h032036: out <= 1'b1;
24'h039036: out <= 1'b1;
24'h03a036: out <= 1'b1;
24'h03b036: out <= 1'b1;
24'h03e036: out <= 1'b1;
24'h03f036: out <= 1'b1;
24'h040036: out <= 1'b1;
24'h04c036: out <= 1'b1;
24'h04d036: out <= 1'b1;
24'h04e036: out <= 1'b1;
24'h04f036: out <= 1'b1;
24'h052036: out <= 1'b1;
24'h053036: out <= 1'b1;
24'h054036: out <= 1'b1;
24'h055036: out <= 1'b1;
24'h056036: out <= 1'b1;
24'h005037: out <= 1'b1;
24'h006037: out <= 1'b1;
24'h010037: out <= 1'b1;
24'h011037: out <= 1'b1;
24'h012037: out <= 1'b1;
24'h01a037: out <= 1'b1;
24'h01b037: out <= 1'b1;
24'h01c037: out <= 1'b1;
24'h021037: out <= 1'b1;
24'h022037: out <= 1'b1;
24'h023037: out <= 1'b1;
24'h024037: out <= 1'b1;
24'h025037: out <= 1'b1;
24'h026037: out <= 1'b1;
24'h027037: out <= 1'b1;
24'h028037: out <= 1'b1;
24'h029037: out <= 1'b1;
24'h030037: out <= 1'b1;
24'h031037: out <= 1'b1;
24'h032037: out <= 1'b1;
24'h033037: out <= 1'b1;
24'h034037: out <= 1'b1;
24'h036037: out <= 1'b1;
24'h037037: out <= 1'b1;
24'h038037: out <= 1'b1;
24'h039037: out <= 1'b1;
24'h03a037: out <= 1'b1;
24'h03b037: out <= 1'b1;
24'h03e037: out <= 1'b1;
24'h03f037: out <= 1'b1;
24'h040037: out <= 1'b1;
24'h041037: out <= 1'b1;
24'h042037: out <= 1'b1;
24'h043037: out <= 1'b1;
24'h044037: out <= 1'b1;
24'h045037: out <= 1'b1;
24'h046037: out <= 1'b1;
24'h047037: out <= 1'b1;
24'h04c037: out <= 1'b1;
24'h04d037: out <= 1'b1;
24'h04e037: out <= 1'b1;
24'h04f037: out <= 1'b1;
24'h050037: out <= 1'b1;
24'h051037: out <= 1'b1;
24'h052037: out <= 1'b1;
24'h053037: out <= 1'b1;
24'h054037: out <= 1'b1;
24'h055037: out <= 1'b1;
24'h005038: out <= 1'b1;
24'h006038: out <= 1'b1;
24'h010038: out <= 1'b1;
24'h011038: out <= 1'b1;
24'h012038: out <= 1'b1;
24'h01b038: out <= 1'b1;
24'h01c038: out <= 1'b1;
24'h023038: out <= 1'b1;
24'h024038: out <= 1'b1;
24'h025038: out <= 1'b1;
24'h026038: out <= 1'b1;
24'h027038: out <= 1'b1;
24'h028038: out <= 1'b1;
24'h030038: out <= 1'b1;
24'h031038: out <= 1'b1;
24'h032038: out <= 1'b1;
24'h033038: out <= 1'b1;
24'h034038: out <= 1'b1;
24'h035038: out <= 1'b1;
24'h036038: out <= 1'b1;
24'h037038: out <= 1'b1;
24'h038038: out <= 1'b1;
24'h039038: out <= 1'b1;
24'h03a038: out <= 1'b1;
24'h03f038: out <= 1'b1;
24'h040038: out <= 1'b1;
24'h041038: out <= 1'b1;
24'h042038: out <= 1'b1;
24'h043038: out <= 1'b1;
24'h044038: out <= 1'b1;
24'h045038: out <= 1'b1;
24'h046038: out <= 1'b1;
24'h047038: out <= 1'b1;
24'h04d038: out <= 1'b1;
24'h04e038: out <= 1'b1;
24'h04f038: out <= 1'b1;
24'h050038: out <= 1'b1;
24'h051038: out <= 1'b1;
24'h052038: out <= 1'b1;
24'h053038: out <= 1'b1;
24'h054038: out <= 1'b1;
24'h031039: out <= 1'b1;
24'h032039: out <= 1'b1;
24'h033039: out <= 1'b1;
24'h034039: out <= 1'b1;
24'h035039: out <= 1'b1;
24'h036039: out <= 1'b1;
24'h037039: out <= 1'b1;
24'h038039: out <= 1'b1;
default: out <= 1'b0;

endcase 
end 
endmodule 